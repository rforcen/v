// assorted collection of polyhedrons
// from https://dmccooey.com/polyhedra/

module poly

pub const depot = [
	Polyhedron{
		name:      'MedialPentagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.7612882
			y: 0.0
			z: 1.231790
		}, Vertex{
			x: 0.7612882
			y: 0.0
			z: -1.231790
		}, Vertex{
			x: -0.7612882
			y: 0.0
			z: 1.231790
		}, Vertex{
			x: -0.7612882
			y: 0.0
			z: -1.231790
		}, Vertex{
			x: 1.231790
			y: 0.7612882
			z: 0.0
		}, Vertex{
			x: 1.231790
			y: -0.7612882
			z: 0.0
		}, Vertex{
			x: -1.231790
			y: 0.7612882
			z: 0.0
		}, Vertex{
			x: -1.231790
			y: -0.7612882
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.231790
			z: 0.7612882
		}, Vertex{
			x: 0.0
			y: 1.231790
			z: -0.7612882
		}, Vertex{
			x: 0.0
			y: -1.231790
			z: 0.7612882
		}, Vertex{
			x: 0.0
			y: -1.231790
			z: -0.7612882
		}, Vertex{
			x: 0.2329835
			y: -0.1855579
			z: 1.172262
		}, Vertex{
			x: 0.2329835
			y: 0.1855579
			z: -1.172262
		}, Vertex{
			x: -0.2329835
			y: 0.1855579
			z: 1.172262
		}, Vertex{
			x: -0.2329835
			y: -0.1855579
			z: -1.172262
		}, Vertex{
			x: 1.172262
			y: -0.2329835
			z: 0.1855579
		}, Vertex{
			x: 1.172262
			y: 0.2329835
			z: -0.1855579
		}, Vertex{
			x: -1.172262
			y: 0.2329835
			z: 0.1855579
		}, Vertex{
			x: -1.172262
			y: -0.2329835
			z: -0.1855579
		}, Vertex{
			x: 0.1855579
			y: -1.172262
			z: 0.2329835
		}, Vertex{
			x: 0.1855579
			y: 1.172262
			z: -0.2329835
		}, Vertex{
			x: -0.1855579
			y: 1.172262
			z: 0.2329835
		}, Vertex{
			x: -0.1855579
			y: -1.172262
			z: -0.2329835
		}, Vertex{
			x: 0.328621
			y: 0.3403026
			z: 1.113154
		}, Vertex{
			x: 0.328621
			y: -0.3403026
			z: -1.113154
		}, Vertex{
			x: -0.328621
			y: -0.3403026
			z: 1.113154
		}, Vertex{
			x: -0.328621
			y: 0.3403026
			z: -1.113154
		}, Vertex{
			x: 1.113154
			y: 0.328621
			z: 0.3403026
		}, Vertex{
			x: 1.113154
			y: -0.328621
			z: -0.3403026
		}, Vertex{
			x: -1.113154
			y: -0.328621
			z: 0.3403026
		}, Vertex{
			x: -1.113154
			y: 0.328621
			z: -0.3403026
		}, Vertex{
			x: 0.3403026
			y: 1.113154
			z: 0.328621
		}, Vertex{
			x: 0.3403026
			y: -1.113154
			z: -0.328621
		}, Vertex{
			x: -0.3403026
			y: -1.113154
			z: 0.328621
		}, Vertex{
			x: -0.3403026
			y: 1.113154
			z: -0.328621
		}, Vertex{
			x: 0.6222993
			y: 0.0
			z: 1.006902
		}, Vertex{
			x: 0.6222993
			y: 0.0
			z: -1.006902
		}, Vertex{
			x: -0.6222993
			y: 0.0
			z: 1.006902
		}, Vertex{
			x: -0.6222993
			y: 0.0
			z: -1.006902
		}, Vertex{
			x: 1.006902
			y: 0.6222993
			z: 0.0
		}, Vertex{
			x: 1.006902
			y: -0.6222993
			z: 0.0
		}, Vertex{
			x: -1.006902
			y: 0.6222993
			z: 0.0
		}, Vertex{
			x: -1.006902
			y: -0.6222993
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.006902
			z: 0.6222993
		}, Vertex{
			x: 0.0
			y: 1.006902
			z: -0.6222993
		}, Vertex{
			x: 0.0
			y: -1.006902
			z: 0.6222993
		}, Vertex{
			x: 0.0
			y: -1.006902
			z: -0.6222993
		}, Vertex{
			x: 0.09563752
			y: -0.7172778
			z: 0.9691625
		}, Vertex{
			x: 0.09563752
			y: 0.7172778
			z: -0.9691625
		}, Vertex{
			x: -0.09563752
			y: 0.7172778
			z: 0.9691625
		}, Vertex{
			x: -0.09563752
			y: -0.7172778
			z: -0.9691625
		}, Vertex{
			x: 0.9691625
			y: -0.09563752
			z: 0.7172778
		}, Vertex{
			x: 0.9691625
			y: 0.09563752
			z: -0.7172778
		}, Vertex{
			x: -0.9691625
			y: 0.09563752
			z: 0.7172778
		}, Vertex{
			x: -0.9691625
			y: -0.09563752
			z: -0.7172778
		}, Vertex{
			x: 0.7172778
			y: -0.9691625
			z: 0.09563752
		}, Vertex{
			x: 0.7172778
			y: 0.9691625
			z: -0.09563752
		}, Vertex{
			x: -0.7172778
			y: 0.9691625
			z: 0.09563752
		}, Vertex{
			x: -0.7172778
			y: -0.9691625
			z: -0.09563752
		}, Vertex{
			x: 0.6288599
			y: -0.4549837
			z: 0.9275964
		}, Vertex{
			x: 0.6288599
			y: 0.4549837
			z: -0.9275964
		}, Vertex{
			x: -0.6288599
			y: 0.4549837
			z: 0.9275964
		}, Vertex{
			x: -0.6288599
			y: -0.4549837
			z: -0.9275964
		}, Vertex{
			x: 0.9275964
			y: -0.6288599
			z: 0.4549837
		}, Vertex{
			x: 0.9275964
			y: 0.6288599
			z: -0.4549837
		}, Vertex{
			x: -0.9275964
			y: 0.6288599
			z: 0.4549837
		}, Vertex{
			x: -0.9275964
			y: -0.6288599
			z: -0.4549837
		}, Vertex{
			x: 0.4549837
			y: -0.9275964
			z: 0.6288599
		}, Vertex{
			x: 0.4549837
			y: 0.9275964
			z: -0.6288599
		}, Vertex{
			x: -0.4549837
			y: 0.9275964
			z: 0.6288599
		}, Vertex{
			x: -0.4549837
			y: -0.9275964
			z: -0.6288599
		}, Vertex{
			x: 0.7836047
			y: 0.3958764
			z: 0.8319589
		}, Vertex{
			x: 0.7836047
			y: -0.3958764
			z: -0.8319589
		}, Vertex{
			x: -0.7836047
			y: -0.3958764
			z: 0.8319589
		}, Vertex{
			x: -0.7836047
			y: 0.3958764
			z: -0.8319589
		}, Vertex{
			x: 0.8319589
			y: 0.7836047
			z: 0.3958764
		}, Vertex{
			x: 0.8319589
			y: -0.7836047
			z: -0.3958764
		}, Vertex{
			x: -0.8319589
			y: -0.7836047
			z: 0.3958764
		}, Vertex{
			x: -0.8319589
			y: 0.7836047
			z: -0.3958764
		}, Vertex{
			x: 0.3958764
			y: 0.8319589
			z: 0.7836047
		}, Vertex{
			x: 0.3958764
			y: -0.8319589
			z: -0.7836047
		}, Vertex{
			x: -0.3958764
			y: -0.8319589
			z: 0.7836047
		}, Vertex{
			x: -0.3958764
			y: 0.8319589
			z: -0.7836047
		}]
		faces:     [[0, 16, 17, 40, 76], [0, 76, 32, 44, 50],
			[0, 50, 62, 38, 26], [0, 26, 82, 46, 68], [0, 68, 56, 41, 16],
			[1, 17, 16, 41, 77], [1, 77, 33, 47, 51], [1, 51, 63, 39, 27],
			[1, 27, 83, 45, 69], [1, 69, 57, 40, 17], [2, 18, 19, 43, 78],
			[2, 78, 34, 46, 48], [2, 48, 60, 36, 24], [2, 24, 80, 44, 70],
			[2, 70, 58, 42, 18], [3, 19, 18, 42, 79], [3, 79, 35, 45, 49],
			[3, 49, 61, 37, 25], [3, 25, 81, 47, 71], [3, 71, 59, 43, 19],
			[4, 21, 22, 44, 80], [4, 80, 24, 36, 52], [4, 52, 64, 41, 29],
			[4, 29, 73, 37, 61], [4, 61, 49, 45, 21], [5, 20, 23, 47, 81],
			[5, 81, 25, 37, 53], [5, 53, 65, 40, 28], [5, 28, 72, 36, 60],
			[5, 60, 48, 46, 20], [6, 22, 21, 45, 83], [6, 83, 27, 39, 55],
			[6, 55, 67, 43, 30], [6, 30, 74, 38, 62], [6, 62, 50, 44, 22],
			[7, 23, 20, 46, 82], [7, 82, 26, 38, 54], [7, 54, 66, 42, 31],
			[7, 31, 75, 39, 63], [7, 63, 51, 47, 23], [8, 14, 12, 36, 72],
			[8, 72, 28, 40, 57], [8, 57, 69, 45, 35], [8, 35, 79, 42, 66],
			[8, 66, 54, 38, 14], [9, 13, 15, 39, 75], [9, 75, 31, 42, 58],
			[9, 58, 70, 44, 32], [9, 32, 76, 40, 65], [9, 65, 53, 37, 13],
			[10, 12, 14, 38, 74], [10, 74, 30, 43, 59], [10, 59, 71, 47, 33],
			[10, 33, 77, 41, 64], [10, 64, 52, 36, 12], [11, 15, 13, 37, 73],
			[11, 73, 29, 41, 56], [11, 56, 68, 46, 34], [11, 34, 78, 43, 67],
			[11, 67, 55, 39, 15]]
	},
	Polyhedron{
		name:      'SmallRhombidodecacron'
		vertexes_: [Vertex{
			x: 1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: 2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 2.236068
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -2.236068
		}, Vertex{
			x: 2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.236068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -2.236068
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: -0.690983
		}]
		faces:     [[0, 14, 5, 26], [0, 36, 10, 28], [0, 24, 2, 20],
			[0, 22, 8, 12], [0, 34, 4, 18], [1, 14, 4, 29], [1, 37, 5, 21],
			[1, 25, 11, 13], [1, 23, 3, 19], [1, 35, 9, 27], [2, 15, 6, 32],
			[2, 38, 8, 30], [2, 18, 0, 22], [2, 20, 10, 12], [2, 40, 7, 24],
			[3, 15, 7, 31], [3, 39, 6, 23], [3, 19, 9, 13], [3, 21, 1, 25],
			[3, 41, 11, 33], [4, 16, 9, 34], [4, 19, 1, 35], [4, 29, 5, 27],
			[4, 28, 0, 14], [4, 18, 8, 26], [5, 17, 10, 37], [5, 20, 0, 36],
			[5, 26, 4, 28], [5, 27, 1, 14], [5, 21, 11, 29], [6, 16, 8, 39],
			[6, 22, 2, 38], [6, 32, 7, 30], [6, 33, 3, 15], [6, 23, 9, 31],
			[7, 17, 11, 40], [7, 25, 3, 41], [7, 31, 6, 33], [7, 30, 2, 15],
			[7, 24, 10, 32], [8, 12, 2, 18], [8, 30, 6, 22], [8, 39, 9, 38],
			[8, 35, 4, 16], [8, 26, 0, 34], [9, 13, 1, 23], [9, 27, 4, 19],
			[9, 34, 8, 35], [9, 38, 6, 16], [9, 31, 3, 39], [10, 12, 0, 24],
			[10, 28, 5, 20], [10, 37, 11, 36], [10, 41, 7, 17],
			[10, 32, 2, 40], [11, 13, 3, 21], [11, 33, 7, 25],
			[11, 40, 10, 41], [11, 36, 5, 17], [11, 29, 1, 37]]
	},
	Polyhedron{
		name:      'SnubDodecahedron(laevo}'
		vertexes_: [Vertex{
			x: 0.3748217
			y: -0.3309210
			z: 2.097054
		}, Vertex{
			x: 0.3748217
			y: 0.3309210
			z: -2.097054
		}, Vertex{
			x: -0.3748217
			y: 0.3309210
			z: 2.097054
		}, Vertex{
			x: -0.3748217
			y: -0.3309210
			z: -2.097054
		}, Vertex{
			x: 2.097054
			y: -0.3748217
			z: 0.3309210
		}, Vertex{
			x: 2.097054
			y: 0.3748217
			z: -0.3309210
		}, Vertex{
			x: -2.097054
			y: 0.3748217
			z: 0.3309210
		}, Vertex{
			x: -2.097054
			y: -0.3748217
			z: -0.3309210
		}, Vertex{
			x: 0.3309210
			y: -2.097054
			z: 0.3748217
		}, Vertex{
			x: 0.3309210
			y: 2.097054
			z: -0.3748217
		}, Vertex{
			x: -0.3309210
			y: 2.097054
			z: 0.3748217
		}, Vertex{
			x: -0.3309210
			y: -2.097054
			z: -0.3748217
		}, Vertex{
			x: 0.5677154
			y: 0.6430296
			z: 1.977839
		}, Vertex{
			x: 0.5677154
			y: -0.6430296
			z: -1.977839
		}, Vertex{
			x: -0.5677154
			y: -0.6430296
			z: 1.977839
		}, Vertex{
			x: -0.5677154
			y: 0.6430296
			z: -1.977839
		}, Vertex{
			x: 1.977839
			y: 0.5677154
			z: 0.6430296
		}, Vertex{
			x: 1.977839
			y: -0.5677154
			z: -0.6430296
		}, Vertex{
			x: -1.977839
			y: -0.5677154
			z: 0.6430296
		}, Vertex{
			x: -1.977839
			y: 0.5677154
			z: -0.6430296
		}, Vertex{
			x: 0.6430296
			y: 1.977839
			z: 0.5677154
		}, Vertex{
			x: 0.6430296
			y: -1.977839
			z: -0.5677154
		}, Vertex{
			x: -0.6430296
			y: -1.977839
			z: 0.5677154
		}, Vertex{
			x: -0.6430296
			y: 1.977839
			z: -0.5677154
		}, Vertex{
			x: 0.1928937
			y: -1.249504
			z: 1.746187
		}, Vertex{
			x: 0.1928937
			y: 1.249504
			z: -1.746187
		}, Vertex{
			x: -0.1928937
			y: 1.249504
			z: 1.746187
		}, Vertex{
			x: -0.1928937
			y: -1.249504
			z: -1.746187
		}, Vertex{
			x: 1.746187
			y: -0.1928937
			z: 1.249504
		}, Vertex{
			x: 1.746187
			y: 0.1928937
			z: -1.249504
		}, Vertex{
			x: -1.746187
			y: 0.1928937
			z: 1.249504
		}, Vertex{
			x: -1.746187
			y: -0.1928937
			z: -1.249504
		}, Vertex{
			x: 1.249504
			y: -1.746187
			z: 0.1928937
		}, Vertex{
			x: 1.249504
			y: 1.746187
			z: -0.1928937
		}, Vertex{
			x: -1.249504
			y: 1.746187
			z: 0.1928937
		}, Vertex{
			x: -1.249504
			y: -1.746187
			z: -0.1928937
		}, Vertex{
			x: 1.103157
			y: -0.8475500
			z: 1.646918
		}, Vertex{
			x: 1.103157
			y: 0.8475500
			z: -1.646918
		}, Vertex{
			x: -1.103157
			y: 0.8475500
			z: 1.646918
		}, Vertex{
			x: -1.103157
			y: -0.8475500
			z: -1.646918
		}, Vertex{
			x: 1.646918
			y: -1.103157
			z: 0.8475500
		}, Vertex{
			x: 1.646918
			y: 1.103157
			z: -0.8475500
		}, Vertex{
			x: -1.646918
			y: 1.103157
			z: 0.8475500
		}, Vertex{
			x: -1.646918
			y: -1.103157
			z: -0.8475500
		}, Vertex{
			x: 0.8475500
			y: -1.646918
			z: 1.103157
		}, Vertex{
			x: 0.8475500
			y: 1.646918
			z: -1.103157
		}, Vertex{
			x: -0.8475500
			y: 1.646918
			z: 1.103157
		}, Vertex{
			x: -0.8475500
			y: -1.646918
			z: -1.103157
		}, Vertex{
			x: 1.415265
			y: 0.7283352
			z: 1.454024
		}, Vertex{
			x: 1.415265
			y: -0.7283352
			z: -1.454024
		}, Vertex{
			x: -1.415265
			y: -0.7283352
			z: 1.454024
		}, Vertex{
			x: -1.415265
			y: 0.7283352
			z: -1.454024
		}, Vertex{
			x: 1.454024
			y: 1.415265
			z: 0.7283352
		}, Vertex{
			x: 1.454024
			y: -1.415265
			z: -0.7283352
		}, Vertex{
			x: -1.454024
			y: -1.415265
			z: 0.7283352
		}, Vertex{
			x: -1.454024
			y: 1.415265
			z: -0.7283352
		}, Vertex{
			x: 0.7283352
			y: 1.454024
			z: 1.415265
		}, Vertex{
			x: 0.7283352
			y: -1.454024
			z: -1.415265
		}, Vertex{
			x: -0.7283352
			y: -1.454024
			z: 1.415265
		}, Vertex{
			x: -0.7283352
			y: 1.454024
			z: -1.415265
		}]
		faces:     [[0, 36, 28, 48, 12], [1, 37, 29, 49, 13],
			[2, 38, 30, 50, 14], [3, 39, 31, 51, 15], [4, 40, 32, 53, 17],
			[5, 41, 33, 52, 16], [6, 42, 34, 55, 19], [7, 43, 35, 54, 18],
			[8, 44, 24, 58, 22], [9, 45, 25, 59, 23], [10, 46, 26, 56, 20],
			[11, 47, 27, 57, 21], [0, 2, 14], [1, 3, 15], [2, 0, 12],
			[3, 1, 13], [4, 5, 16], [5, 4, 17], [6, 7, 18], [7, 6, 19],
			[8, 11, 21], [9, 10, 20], [10, 9, 23], [11, 8, 22],
			[12, 48, 56], [13, 49, 57], [14, 50, 58], [15, 51, 59],
			[16, 52, 48], [17, 53, 49], [18, 54, 50], [19, 55, 51],
			[20, 56, 52], [21, 57, 53], [22, 58, 54], [23, 59, 55],
			[24, 44, 36], [25, 45, 37], [26, 46, 38], [27, 47, 39],
			[28, 36, 40], [29, 37, 41], [30, 38, 42], [31, 39, 43],
			[32, 40, 44], [33, 41, 45], [34, 42, 46], [35, 43, 47],
			[36, 0, 24], [37, 1, 25], [38, 2, 26], [39, 3, 27],
			[40, 4, 28], [41, 5, 29], [42, 6, 30], [43, 7, 31],
			[44, 8, 32], [45, 9, 33], [46, 10, 34], [47, 11, 35],
			[48, 28, 16], [49, 29, 17], [50, 30, 18], [51, 31, 19],
			[52, 33, 20], [53, 32, 21], [54, 35, 22], [55, 34, 23],
			[56, 26, 12], [57, 27, 13], [58, 24, 14], [59, 25, 15],
			[24, 0, 14], [25, 1, 15], [26, 2, 12], [27, 3, 13],
			[28, 4, 16], [29, 5, 17], [30, 6, 18], [31, 7, 19],
			[32, 8, 21], [33, 9, 20], [34, 10, 23], [35, 11, 22],
			[36, 44, 40], [37, 45, 41], [38, 46, 42], [39, 47, 43],
			[48, 52, 56], [49, 53, 57], [50, 54, 58], [51, 55, 59]]
	},
	Polyhedron{
		name:      'PentakisDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: 0.927051
			z: -2.427051
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: -2.427051
		}, Vertex{
			x: 2.427051
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: 2.427051
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: 0.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: 0.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: 1.330587
			y: 0.0
			z: 2.152935
		}, Vertex{
			x: 1.330587
			y: 0.0
			z: -2.152935
		}, Vertex{
			x: -1.330587
			y: 0.0
			z: 2.152935
		}, Vertex{
			x: -1.330587
			y: 0.0
			z: -2.152935
		}, Vertex{
			x: 2.152935
			y: 1.330587
			z: 0.0
		}, Vertex{
			x: 2.152935
			y: -1.330587
			z: 0.0
		}, Vertex{
			x: -2.152935
			y: 1.330587
			z: 0.0
		}, Vertex{
			x: -2.152935
			y: -1.330587
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.152935
			z: 1.330587
		}, Vertex{
			x: 0.0
			y: 2.152935
			z: -1.330587
		}, Vertex{
			x: 0.0
			y: -2.152935
			z: 1.330587
		}, Vertex{
			x: 0.0
			y: -2.152935
			z: -1.330587
		}, Vertex{
			x: 1.5
			y: 1.5
			z: 1.5
		}, Vertex{
			x: 1.5
			y: 1.5
			z: -1.5
		}, Vertex{
			x: 1.5
			y: -1.5
			z: 1.5
		}, Vertex{
			x: 1.5
			y: -1.5
			z: -1.5
		}, Vertex{
			x: -1.5
			y: 1.5
			z: 1.5
		}, Vertex{
			x: -1.5
			y: 1.5
			z: -1.5
		}, Vertex{
			x: -1.5
			y: -1.5
			z: 1.5
		}, Vertex{
			x: -1.5
			y: -1.5
			z: -1.5
		}]
		faces:     [[12, 0, 2], [12, 2, 26], [12, 26, 4], [12, 4, 24],
			[12, 24, 0], [13, 3, 1], [13, 1, 25], [13, 25, 5],
			[13, 5, 27], [13, 27, 3], [14, 2, 0], [14, 0, 28],
			[14, 28, 6], [14, 6, 30], [14, 30, 2], [15, 1, 3],
			[15, 3, 31], [15, 31, 7], [15, 7, 29], [15, 29, 1],
			[16, 4, 5], [16, 5, 25], [16, 25, 8], [16, 8, 24],
			[16, 24, 4], [17, 5, 4], [17, 4, 26], [17, 26, 9],
			[17, 9, 27], [17, 27, 5], [18, 7, 6], [18, 6, 28],
			[18, 28, 10], [18, 10, 29], [18, 29, 7], [19, 6, 7],
			[19, 7, 31], [19, 31, 11], [19, 11, 30], [19, 30, 6],
			[20, 8, 10], [20, 10, 28], [20, 28, 0], [20, 0, 24],
			[20, 24, 8], [21, 10, 8], [21, 8, 25], [21, 25, 1],
			[21, 1, 29], [21, 29, 10], [22, 11, 9], [22, 9, 26],
			[22, 26, 2], [22, 2, 30], [22, 30, 11], [23, 9, 11],
			[23, 11, 31], [23, 31, 3], [23, 3, 27], [23, 27, 9]]
	},
	Polyhedron{
		name:      'SmallSnubIcosicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.2678437
			y: 0.0
			z: 1.433380
		}, Vertex{
			x: 0.2678437
			y: 0.0
			z: -1.433380
		}, Vertex{
			x: -0.2678437
			y: 0.0
			z: 1.433380
		}, Vertex{
			x: -0.2678437
			y: 0.0
			z: -1.433380
		}, Vertex{
			x: 1.433380
			y: 0.2678437
			z: 0.0
		}, Vertex{
			x: 1.433380
			y: -0.2678437
			z: 0.0
		}, Vertex{
			x: -1.433380
			y: 0.2678437
			z: 0.0
		}, Vertex{
			x: -1.433380
			y: -0.2678437
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.433380
			z: 0.2678437
		}, Vertex{
			x: 0.0
			y: 1.433380
			z: -0.2678437
		}, Vertex{
			x: 0.0
			y: -1.433380
			z: 0.2678437
		}, Vertex{
			x: 0.0
			y: -1.433380
			z: -0.2678437
		}, Vertex{
			x: 0.5768607
			y: 0.5
			z: 1.242397
		}, Vertex{
			x: 0.5768607
			y: 0.5
			z: -1.242397
		}, Vertex{
			x: 0.5768607
			y: -0.5
			z: 1.242397
		}, Vertex{
			x: 0.5768607
			y: -0.5
			z: -1.242397
		}, Vertex{
			x: -0.5768607
			y: 0.5
			z: 1.242397
		}, Vertex{
			x: -0.5768607
			y: 0.5
			z: -1.242397
		}, Vertex{
			x: -0.5768607
			y: -0.5
			z: 1.242397
		}, Vertex{
			x: -0.5768607
			y: -0.5
			z: -1.242397
		}, Vertex{
			x: 1.242397
			y: 0.5768607
			z: 0.5
		}, Vertex{
			x: 1.242397
			y: 0.5768607
			z: -0.5
		}, Vertex{
			x: 1.242397
			y: -0.5768607
			z: 0.5
		}, Vertex{
			x: 1.242397
			y: -0.5768607
			z: -0.5
		}, Vertex{
			x: -1.242397
			y: 0.5768607
			z: 0.5
		}, Vertex{
			x: -1.242397
			y: 0.5768607
			z: -0.5
		}, Vertex{
			x: -1.242397
			y: -0.5768607
			z: 0.5
		}, Vertex{
			x: -1.242397
			y: -0.5768607
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.242397
			z: 0.5768607
		}, Vertex{
			x: 0.5
			y: 1.242397
			z: -0.5768607
		}, Vertex{
			x: 0.5
			y: -1.242397
			z: 0.5768607
		}, Vertex{
			x: 0.5
			y: -1.242397
			z: -0.5768607
		}, Vertex{
			x: -0.5
			y: 1.242397
			z: 0.5768607
		}, Vertex{
			x: -0.5
			y: 1.242397
			z: -0.5768607
		}, Vertex{
			x: -0.5
			y: -1.242397
			z: 0.5768607
		}, Vertex{
			x: -0.5
			y: -1.242397
			z: -0.5768607
		}, Vertex{
			x: 0.309017
			y: 0.9333802
			z: 1.076861
		}, Vertex{
			x: 0.309017
			y: 0.9333802
			z: -1.076861
		}, Vertex{
			x: 0.309017
			y: -0.9333802
			z: 1.076861
		}, Vertex{
			x: 0.309017
			y: -0.9333802
			z: -1.076861
		}, Vertex{
			x: -0.309017
			y: 0.9333802
			z: 1.076861
		}, Vertex{
			x: -0.309017
			y: 0.9333802
			z: -1.076861
		}, Vertex{
			x: -0.309017
			y: -0.9333802
			z: 1.076861
		}, Vertex{
			x: -0.309017
			y: -0.9333802
			z: -1.076861
		}, Vertex{
			x: 1.076861
			y: 0.309017
			z: 0.9333802
		}, Vertex{
			x: 1.076861
			y: 0.309017
			z: -0.9333802
		}, Vertex{
			x: 1.076861
			y: -0.309017
			z: 0.9333802
		}, Vertex{
			x: 1.076861
			y: -0.309017
			z: -0.9333802
		}, Vertex{
			x: -1.076861
			y: 0.309017
			z: 0.9333802
		}, Vertex{
			x: -1.076861
			y: 0.309017
			z: -0.9333802
		}, Vertex{
			x: -1.076861
			y: -0.309017
			z: 0.9333802
		}, Vertex{
			x: -1.076861
			y: -0.309017
			z: -0.9333802
		}, Vertex{
			x: 0.9333802
			y: 1.076861
			z: 0.309017
		}, Vertex{
			x: 0.9333802
			y: 1.076861
			z: -0.309017
		}, Vertex{
			x: 0.9333802
			y: -1.076861
			z: 0.309017
		}, Vertex{
			x: 0.9333802
			y: -1.076861
			z: -0.309017
		}, Vertex{
			x: -0.9333802
			y: 1.076861
			z: 0.309017
		}, Vertex{
			x: -0.9333802
			y: 1.076861
			z: -0.309017
		}, Vertex{
			x: -0.9333802
			y: -1.076861
			z: 0.309017
		}, Vertex{
			x: -0.9333802
			y: -1.076861
			z: -0.309017
		}]
		faces:     [[0, 46, 12, 14, 44], [1, 45, 15, 13, 47],
			[2, 48, 18, 16, 50], [3, 51, 17, 19, 49], [4, 53, 20, 21, 52],
			[5, 54, 23, 22, 55], [6, 56, 25, 24, 57], [7, 59, 26, 27, 58],
			[8, 40, 28, 32, 36], [9, 37, 33, 29, 41], [10, 38, 34, 30, 42],
			[11, 43, 31, 35, 39], [0, 16, 18], [1, 19, 17], [2, 14, 12],
			[3, 13, 15], [4, 22, 23], [5, 21, 20], [6, 27, 26],
			[7, 24, 25], [8, 29, 33], [9, 32, 28], [10, 35, 31],
			[11, 30, 34], [12, 28, 40], [13, 41, 29], [14, 42, 30],
			[15, 31, 43], [16, 36, 32], [17, 33, 37], [18, 34, 38],
			[19, 39, 35], [20, 12, 46], [21, 47, 13], [22, 44, 14],
			[23, 15, 45], [24, 50, 16], [25, 17, 51], [26, 18, 48],
			[27, 49, 19], [28, 20, 53], [29, 52, 21], [30, 55, 22],
			[31, 23, 54], [32, 57, 24], [33, 25, 56], [34, 26, 59],
			[35, 58, 27], [36, 0, 44], [37, 45, 1], [38, 46, 0],
			[39, 1, 47], [40, 48, 2], [41, 3, 49], [42, 2, 50],
			[43, 51, 3], [44, 4, 52], [45, 53, 4], [46, 54, 5],
			[47, 5, 55], [48, 56, 6], [49, 6, 57], [50, 7, 58],
			[51, 59, 7], [52, 8, 36], [53, 37, 9], [54, 38, 10],
			[55, 11, 39], [56, 40, 8], [57, 9, 41], [58, 10, 42],
			[59, 43, 11], [0, 18, 38], [0, 36, 16], [1, 17, 37],
			[1, 39, 19], [2, 12, 40], [2, 42, 14], [3, 15, 43],
			[3, 41, 13], [21, 5, 47], [21, 13, 29], [22, 4, 44],
			[22, 14, 30], [25, 33, 17], [25, 51, 7], [26, 34, 18],
			[26, 48, 6], [28, 12, 20], [28, 53, 9], [31, 15, 23],
			[31, 54, 10], [32, 9, 57], [32, 24, 16], [35, 10, 58],
			[35, 27, 19], [45, 4, 23], [45, 37, 53], [46, 5, 20],
			[46, 38, 54], [49, 27, 6], [49, 57, 41], [50, 24, 7],
			[50, 58, 42], [52, 29, 8], [52, 36, 44], [55, 30, 11],
			[55, 39, 47], [56, 8, 33], [56, 48, 40], [59, 11, 34],
			[59, 51, 43]]
	},
	Polyhedron{
		name:      'Rhombicuboctahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: -0.5
		}]
		faces:     [[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9],
			[12, 13, 15, 14], [16, 17, 21, 20], [18, 22, 23, 19],
			[0, 2, 10, 8], [0, 16, 20, 4], [7, 3, 19, 23], [7, 15, 13, 5],
			[11, 3, 1, 9], [11, 10, 18, 19], [12, 14, 6, 4], [12, 20, 21, 13],
			[17, 1, 5, 21], [17, 16, 8, 9], [22, 14, 15, 23],
			[22, 18, 2, 6], [0, 8, 16], [1, 17, 9], [2, 18, 10],
			[3, 11, 19], [4, 20, 12], [5, 13, 21], [6, 14, 22],
			[7, 23, 15]]
	},
	Polyhedron{
		name:      'GreatPentagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.2163811
			y: -0.2395588
			z: 0.6449711
		}, Vertex{
			x: -0.2163811
			y: -0.2395588
			z: -0.6449711
		}, Vertex{
			x: -0.2163811
			y: 0.2395588
			z: 0.6449711
		}, Vertex{
			x: 0.2163811
			y: 0.2395588
			z: -0.6449711
		}, Vertex{
			x: -0.2395588
			y: 0.6449711
			z: 0.2163811
		}, Vertex{
			x: 0.2395588
			y: 0.6449711
			z: -0.2163811
		}, Vertex{
			x: 0.2395588
			y: -0.6449711
			z: 0.2163811
		}, Vertex{
			x: -0.2395588
			y: -0.6449711
			z: -0.2163811
		}, Vertex{
			x: 0.6449711
			y: 0.2163811
			z: -0.2395588
		}, Vertex{
			x: -0.6449711
			y: 0.2163811
			z: 0.2395588
		}, Vertex{
			x: -0.6449711
			y: -0.2163811
			z: -0.2395588
		}, Vertex{
			x: 0.6449711
			y: -0.2163811
			z: 0.2395588
		}, Vertex{
			x: 0.6737688
			y: 0.0
			z: 0.2573568
		}, Vertex{
			x: 0.6737688
			y: 0.0
			z: -0.2573568
		}, Vertex{
			x: -0.6737688
			y: 0.0
			z: 0.2573568
		}, Vertex{
			x: -0.6737688
			y: 0.0
			z: -0.2573568
		}, Vertex{
			x: 0.0
			y: 0.2573568
			z: 0.6737688
		}, Vertex{
			x: 0.0
			y: 0.2573568
			z: -0.6737688
		}, Vertex{
			x: 0.0
			y: -0.2573568
			z: 0.6737688
		}, Vertex{
			x: 0.0
			y: -0.2573568
			z: -0.6737688
		}, Vertex{
			x: 0.2573568
			y: 0.6737688
			z: 0.0
		}, Vertex{
			x: -0.2573568
			y: 0.6737688
			z: 0.0
		}, Vertex{
			x: 0.2573568
			y: -0.6737688
			z: 0.0
		}, Vertex{
			x: -0.2573568
			y: -0.6737688
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.5669247
			z: 0.3503788
		}, Vertex{
			x: 0.0
			y: -0.5669247
			z: -0.3503788
		}, Vertex{
			x: 0.0
			y: 0.5669247
			z: 0.3503788
		}, Vertex{
			x: 0.0
			y: 0.5669247
			z: -0.3503788
		}, Vertex{
			x: -0.5669247
			y: 0.3503788
			z: 0.0
		}, Vertex{
			x: 0.5669247
			y: 0.3503788
			z: 0.0
		}, Vertex{
			x: -0.5669247
			y: -0.3503788
			z: 0.0
		}, Vertex{
			x: 0.5669247
			y: -0.3503788
			z: 0.0
		}, Vertex{
			x: 0.3503788
			y: 0.0
			z: -0.5669247
		}, Vertex{
			x: 0.3503788
			y: 0.0
			z: 0.5669247
		}, Vertex{
			x: -0.3503788
			y: 0.0
			z: -0.5669247
		}, Vertex{
			x: -0.3503788
			y: 0.0
			z: 0.5669247
		}, Vertex{
			x: -0.4235137
			y: -0.5747065
			z: 0.1026907
		}, Vertex{
			x: 0.4235137
			y: -0.5747065
			z: -0.1026907
		}, Vertex{
			x: 0.4235137
			y: 0.5747065
			z: 0.1026907
		}, Vertex{
			x: -0.4235137
			y: 0.5747065
			z: -0.1026907
		}, Vertex{
			x: 0.5747065
			y: 0.1026907
			z: 0.4235137
		}, Vertex{
			x: -0.5747065
			y: 0.1026907
			z: -0.4235137
		}, Vertex{
			x: -0.5747065
			y: -0.1026907
			z: 0.4235137
		}, Vertex{
			x: 0.5747065
			y: -0.1026907
			z: -0.4235137
		}, Vertex{
			x: -0.1026907
			y: 0.4235137
			z: -0.5747065
		}, Vertex{
			x: 0.1026907
			y: 0.4235137
			z: 0.5747065
		}, Vertex{
			x: 0.1026907
			y: -0.4235137
			z: -0.5747065
		}, Vertex{
			x: -0.1026907
			y: -0.4235137
			z: 0.5747065
		}, Vertex{
			x: 0.5715693
			y: -0.3351477
			z: -0.2849236
		}, Vertex{
			x: -0.5715693
			y: -0.3351477
			z: 0.2849236
		}, Vertex{
			x: -0.5715693
			y: 0.3351477
			z: -0.2849236
		}, Vertex{
			x: 0.5715693
			y: 0.3351477
			z: 0.2849236
		}, Vertex{
			x: -0.3351477
			y: -0.2849236
			z: 0.5715693
		}, Vertex{
			x: 0.3351477
			y: -0.2849236
			z: -0.5715693
		}, Vertex{
			x: 0.3351477
			y: 0.2849236
			z: 0.5715693
		}, Vertex{
			x: -0.3351477
			y: 0.2849236
			z: -0.5715693
		}, Vertex{
			x: -0.2849236
			y: 0.5715693
			z: -0.3351477
		}, Vertex{
			x: 0.2849236
			y: 0.5715693
			z: 0.3351477
		}, Vertex{
			x: 0.2849236
			y: -0.5715693
			z: -0.3351477
		}, Vertex{
			x: -0.2849236
			y: -0.5715693
			z: 0.3351477
		}, Vertex{
			x: 0.07340182
			y: -0.7084374
			z: -0.1136904
		}, Vertex{
			x: -0.07340182
			y: -0.7084374
			z: 0.1136904
		}, Vertex{
			x: -0.07340182
			y: 0.7084374
			z: -0.1136904
		}, Vertex{
			x: 0.07340182
			y: 0.7084374
			z: 0.1136904
		}, Vertex{
			x: -0.7084374
			y: -0.1136904
			z: 0.07340182
		}, Vertex{
			x: 0.7084374
			y: -0.1136904
			z: -0.07340182
		}, Vertex{
			x: 0.7084374
			y: 0.1136904
			z: 0.07340182
		}, Vertex{
			x: -0.7084374
			y: 0.1136904
			z: -0.07340182
		}, Vertex{
			x: -0.1136904
			y: 0.07340182
			z: -0.7084374
		}, Vertex{
			x: 0.1136904
			y: 0.07340182
			z: 0.7084374
		}, Vertex{
			x: 0.1136904
			y: -0.07340182
			z: -0.7084374
		}, Vertex{
			x: -0.1136904
			y: -0.07340182
			z: 0.7084374
		}, Vertex{
			x: -0.2214573
			y: -0.4688786
			z: -0.5013047
		}, Vertex{
			x: 0.2214573
			y: -0.4688786
			z: 0.5013047
		}, Vertex{
			x: 0.2214573
			y: 0.4688786
			z: -0.5013047
		}, Vertex{
			x: -0.2214573
			y: 0.4688786
			z: 0.5013047
		}, Vertex{
			x: 0.4688786
			y: -0.5013047
			z: 0.2214573
		}, Vertex{
			x: -0.4688786
			y: -0.5013047
			z: -0.2214573
		}, Vertex{
			x: -0.4688786
			y: 0.5013047
			z: 0.2214573
		}, Vertex{
			x: 0.4688786
			y: 0.5013047
			z: -0.2214573
		}, Vertex{
			x: 0.5013047
			y: 0.2214573
			z: -0.4688786
		}, Vertex{
			x: -0.5013047
			y: 0.2214573
			z: 0.4688786
		}, Vertex{
			x: -0.5013047
			y: -0.2214573
			z: -0.4688786
		}, Vertex{
			x: 0.5013047
			y: -0.2214573
			z: 0.4688786
		}, Vertex{
			x: -0.416412
			y: -0.416412
			z: -0.416412
		}, Vertex{
			x: -0.416412
			y: -0.416412
			z: 0.416412
		}, Vertex{
			x: 0.416412
			y: -0.416412
			z: -0.416412
		}, Vertex{
			x: 0.416412
			y: -0.416412
			z: 0.416412
		}, Vertex{
			x: -0.416412
			y: 0.416412
			z: -0.416412
		}, Vertex{
			x: -0.416412
			y: 0.416412
			z: 0.416412
		}, Vertex{
			x: 0.416412
			y: 0.416412
			z: -0.416412
		}, Vertex{
			x: 0.416412
			y: 0.416412
			z: 0.416412
		}]
		faces:     [[24, 0, 2, 14, 36], [24, 36, 72, 86, 76],
			[24, 76, 40, 16, 52], [24, 52, 64, 84, 60], [24, 60, 48, 12, 0],
			[25, 1, 3, 13, 37], [25, 37, 73, 85, 77], [25, 77, 41, 17, 53],
			[25, 53, 65, 87, 61], [25, 61, 49, 15, 1], [26, 2, 0, 12, 38],
			[26, 38, 74, 88, 78], [26, 78, 42, 18, 54], [26, 54, 66, 90, 62],
			[26, 62, 50, 14, 2], [27, 3, 1, 15, 39], [27, 39, 75, 91, 79],
			[27, 79, 43, 19, 55], [27, 55, 67, 89, 63], [27, 63, 51, 13, 3],
			[28, 4, 5, 17, 41], [28, 41, 77, 85, 81], [28, 81, 45, 20, 56],
			[28, 56, 68, 84, 64], [28, 64, 52, 16, 4], [29, 5, 4, 16, 40],
			[29, 40, 76, 86, 80], [29, 80, 44, 21, 57], [29, 57, 69, 87, 65],
			[29, 65, 53, 17, 5], [30, 7, 6, 18, 42], [30, 42, 78, 88, 82],
			[30, 82, 46, 22, 59], [30, 59, 71, 89, 67], [30, 67, 55, 19, 7],
			[31, 6, 7, 19, 43], [31, 43, 79, 91, 83], [31, 83, 47, 23, 58],
			[31, 58, 70, 90, 66], [31, 66, 54, 18, 6], [32, 8, 11, 22, 46],
			[32, 46, 82, 88, 74], [32, 74, 38, 12, 48], [32, 48, 60, 84, 68],
			[32, 68, 56, 20, 8], [33, 11, 8, 20, 45], [33, 45, 81, 85, 73],
			[33, 73, 37, 13, 51], [33, 51, 63, 89, 71], [33, 71, 59, 22, 11],
			[34, 10, 9, 21, 44], [34, 44, 80, 86, 72], [34, 72, 36, 14, 50],
			[34, 50, 62, 90, 70], [34, 70, 58, 23, 10], [35, 9, 10, 23, 47],
			[35, 47, 83, 91, 75], [35, 75, 39, 15, 49], [35, 49, 61, 87, 69],
			[35, 69, 57, 21, 9]]
	},
	Polyhedron{
		name:      'GreatRhombidodecahedron'
		vertexes_: [Vertex{
			x: -0.5
			y: -0.5
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 0.1909830
		}, Vertex{
			x: -0.690983
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: 0.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: -0.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: 0.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.1909830
			y: 0.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: 0.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: 0.618034
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: -0.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: -0.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: -0.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: -0.618034
			z: -0.309017
		}, Vertex{
			x: 0.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: -0.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: -0.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: 0.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.618034
			y: -0.309017
			z: 0.1909830
		}, Vertex{
			x: -0.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: -0.618034
			y: -0.309017
			z: 0.1909830
		}]
		faces:     [[0, 24, 56, 48, 12, 14, 50, 58, 26, 2], [0, 36, 44, 32, 17, 21, 34, 48, 40,
			4],
			[7, 3, 39, 47, 33, 18, 22, 35, 51, 43], [7, 5, 25, 53, 45, 9, 11, 47, 55, 27],
			[10, 8, 44, 52, 24, 4, 6, 26, 54, 46], [10, 11, 29, 37, 53, 17, 16, 52, 36, 28],
			[13, 31, 43, 59, 23, 22, 58, 42, 30, 12], [13, 49, 57, 25, 1, 3, 27, 59, 51, 15],
			[19, 33, 46, 38, 2, 6, 42, 50, 35, 23], [19, 55, 39, 29, 9, 8, 28, 38, 54, 18],
			[20, 16, 32, 45, 37, 1, 5, 41, 49, 34], [20, 21, 57, 41, 31, 15, 14, 30, 40, 56],
			[24, 0, 36, 52], [24, 56, 40, 4], [25, 5, 41, 57],
			[25, 53, 37, 1], [26, 6, 42, 58], [26, 54, 38, 2],
			[27, 3, 39, 55], [27, 59, 43, 7], [28, 8, 44, 36],
			[28, 38, 46, 10], [29, 11, 47, 39], [29, 37, 45, 9],
			[30, 14, 50, 42], [30, 40, 48, 12], [31, 13, 49, 41],
			[31, 43, 51, 15], [32, 16, 52, 44], [32, 45, 53, 17],
			[33, 19, 55, 47], [33, 46, 54, 18], [34, 21, 57, 49],
			[34, 48, 56, 20], [35, 22, 58, 50], [35, 51, 59, 23],
			[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9], [12, 13, 15, 14],
			[16, 17, 21, 20], [18, 22, 23, 19]]
	},
	Polyhedron{
		name:      'Cubohemioctahedron'
		vertexes_: [Vertex{
			x: 0.7071068
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: 0.7071068
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: -0.7071068
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: -0.7071068
		}]
		faces:     [[0, 4, 9, 3, 7, 10], [0, 5, 11, 3, 6, 8],
			[1, 4, 8, 2, 7, 11], [1, 5, 10, 2, 6, 9], [0, 5, 1, 4],
			[0, 8, 2, 10], [7, 2, 6, 3], [7, 11, 5, 10], [9, 1, 11, 3],
			[9, 6, 8, 4]]
	},
	Polyhedron{
		name:      'GreatStellapentakisDodecahedron'
		vertexes_: [Vertex{
			x: 2.427051
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: 2.427051
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: 0.0
			y: 0.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: 0.927051
			z: -2.427051
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: -2.427051
		}, Vertex{
			x: 0.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: 0.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.8009920
			z: 0.4950402
		}, Vertex{
			x: 0.0
			y: -0.8009920
			z: -0.4950402
		}, Vertex{
			x: 0.0
			y: 0.8009920
			z: 0.4950402
		}, Vertex{
			x: 0.0
			y: 0.8009920
			z: -0.4950402
		}, Vertex{
			x: -0.8009920
			y: 0.4950402
			z: 0.0
		}, Vertex{
			x: 0.8009920
			y: 0.4950402
			z: 0.0
		}, Vertex{
			x: -0.8009920
			y: -0.4950402
			z: 0.0
		}, Vertex{
			x: 0.8009920
			y: -0.4950402
			z: 0.0
		}, Vertex{
			x: 0.4950402
			y: 0.0
			z: -0.8009920
		}, Vertex{
			x: 0.4950402
			y: 0.0
			z: 0.8009920
		}, Vertex{
			x: -0.4950402
			y: 0.0
			z: -0.8009920
		}, Vertex{
			x: -0.4950402
			y: 0.0
			z: 0.8009920
		}, Vertex{
			x: -1.5
			y: -1.5
			z: -1.5
		}, Vertex{
			x: -1.5
			y: -1.5
			z: 1.5
		}, Vertex{
			x: 1.5
			y: -1.5
			z: -1.5
		}, Vertex{
			x: 1.5
			y: -1.5
			z: 1.5
		}, Vertex{
			x: -1.5
			y: 1.5
			z: -1.5
		}, Vertex{
			x: -1.5
			y: 1.5
			z: 1.5
		}, Vertex{
			x: 1.5
			y: 1.5
			z: -1.5
		}, Vertex{
			x: 1.5
			y: 1.5
			z: 1.5
		}]
		faces:     [[12, 0, 2], [12, 2, 26], [12, 26, 4], [12, 4, 24],
			[12, 24, 0], [13, 3, 1], [13, 1, 25], [13, 25, 5],
			[13, 5, 27], [13, 27, 3], [14, 2, 0], [14, 0, 28],
			[14, 28, 6], [14, 6, 30], [14, 30, 2], [15, 1, 3],
			[15, 3, 31], [15, 31, 7], [15, 7, 29], [15, 29, 1],
			[16, 4, 5], [16, 5, 25], [16, 25, 8], [16, 8, 24],
			[16, 24, 4], [17, 5, 4], [17, 4, 26], [17, 26, 9],
			[17, 9, 27], [17, 27, 5], [18, 7, 6], [18, 6, 28],
			[18, 28, 10], [18, 10, 29], [18, 29, 7], [19, 6, 7],
			[19, 7, 31], [19, 31, 11], [19, 11, 30], [19, 30, 6],
			[20, 8, 10], [20, 10, 28], [20, 28, 0], [20, 0, 24],
			[20, 24, 8], [21, 10, 8], [21, 8, 25], [21, 25, 1],
			[21, 1, 29], [21, 29, 10], [22, 11, 9], [22, 9, 26],
			[22, 26, 2], [22, 2, 30], [22, 30, 11], [23, 9, 11],
			[23, 11, 31], [23, 31, 3], [23, 3, 27], [23, 27, 9]]
	},
	Polyhedron{
		name:      'UniformGreatRhombicuboctahedron'
		vertexes_: [Vertex{
			x: -0.5
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: 0.5
		}]
		faces:     [[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9],
			[12, 13, 15, 14], [16, 17, 21, 20], [18, 22, 23, 19],
			[0, 2, 10, 8], [0, 16, 20, 4], [7, 3, 19, 23], [7, 15, 13, 5],
			[11, 3, 1, 9], [11, 10, 18, 19], [12, 14, 6, 4], [12, 20, 21, 13],
			[17, 1, 5, 21], [17, 16, 8, 9], [22, 14, 15, 23],
			[22, 18, 2, 6], [0, 8, 16], [1, 17, 9], [2, 18, 10],
			[3, 11, 19], [4, 20, 12], [5, 13, 21], [6, 14, 22],
			[7, 23, 15]]
	},
	Polyhedron{
		name:      'GreatTruncatedCuboctahedron'
		vertexes_: [Vertex{
			x: -0.2071068
			y: 0.5
			z: -0.9142135
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: 0.9142135
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: -0.9142135
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: 0.9142135
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: -0.9142135
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: 0.9142135
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: -0.9142135
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: 0.9142135
		}, Vertex{
			x: -0.9142135
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: -0.9142135
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: -0.9142135
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: -0.9142135
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.9142135
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: 0.9142135
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: 0.9142135
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: 0.9142135
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.9142135
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: -0.9142135
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: 0.9142135
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: 0.9142135
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: -0.9142135
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: -0.9142135
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: 0.9142135
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: 0.9142135
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: -0.9142135
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: 0.9142135
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: -0.9142135
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: 0.9142135
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: -0.9142135
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: 0.9142135
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: -0.9142135
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: 0.9142135
		}, Vertex{
			x: -0.9142135
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: -0.9142135
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: -0.9142135
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: -0.9142135
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: 0.9142135
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.9142135
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: 0.9142135
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: 0.9142135
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: -0.2071068
			y: -0.9142135
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: -0.9142135
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: 0.9142135
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: 0.9142135
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: -0.9142135
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: -0.9142135
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: 0.9142135
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: 0.9142135
			z: -0.5
		}]
		faces:     [[0, 24, 28, 4, 6, 30, 26, 2], [1, 3, 27, 31, 7, 5, 29, 25],
			[8, 32, 34, 10, 11, 35, 33, 9], [12, 13, 37, 39, 15, 14, 38, 36],
			[16, 40, 41, 17, 21, 45, 44, 20], [18, 22, 46, 47, 23, 19, 43, 42],
			[0, 32, 8, 40, 16, 24], [1, 25, 17, 41, 9, 33], [2, 26, 18, 42, 10, 34],
			[3, 35, 11, 43, 19, 27], [4, 28, 20, 44, 12, 36],
			[5, 37, 13, 45, 21, 29], [6, 38, 14, 46, 22, 30],
			[7, 31, 23, 47, 15, 39], [0, 2, 34, 32], [1, 33, 35, 3],
			[4, 36, 38, 6], [5, 7, 39, 37], [8, 9, 41, 40], [10, 42, 43, 11],
			[12, 44, 45, 13], [14, 15, 47, 46], [16, 20, 28, 24],
			[17, 25, 29, 21], [18, 26, 30, 22], [19, 23, 31, 27]]
	},
	Polyhedron{
		name:      'SmallDodecicosacron'
		vertexes_: [Vertex{
			x: 2.427051
			y: 0.0
			z: 3.927051
		}, Vertex{
			x: 2.427051
			y: 0.0
			z: -3.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: 3.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: -3.927051
		}, Vertex{
			x: 3.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: 3.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: -3.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: -3.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 3.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: 3.927051
			z: -2.427051
		}, Vertex{
			x: 0.0
			y: -3.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: -3.927051
			z: -2.427051
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: -1.118034
		}]
		faces:     [[0, 18, 6, 14], [0, 22, 9, 12], [0, 25, 1, 24],
			[0, 27, 11, 16], [0, 23, 7, 26], [1, 19, 7, 13], [1, 23, 10, 15],
			[1, 26, 0, 27], [1, 24, 8, 17], [1, 22, 6, 25], [2, 16, 5, 12],
			[2, 21, 11, 14], [2, 31, 3, 30], [2, 29, 9, 18], [2, 20, 4, 28],
			[3, 17, 4, 15], [3, 20, 8, 13], [3, 28, 2, 29], [3, 30, 10, 19],
			[3, 21, 5, 31], [4, 14, 2, 16], [4, 28, 6, 24], [4, 29, 3, 20],
			[4, 15, 11, 25], [4, 21, 10, 17], [5, 12, 8, 26],
			[5, 20, 9, 16], [5, 13, 3, 17], [5, 31, 7, 27], [5, 30, 2, 21],
			[6, 14, 10, 28], [6, 23, 11, 18], [6, 15, 1, 19],
			[6, 25, 4, 29], [6, 24, 0, 22], [7, 12, 0, 18], [7, 26, 5, 30],
			[7, 27, 1, 23], [7, 13, 9, 31], [7, 22, 8, 19], [8, 13, 1, 22],
			[8, 17, 5, 20], [8, 26, 10, 24], [8, 30, 7, 12], [8, 19, 3, 28],
			[9, 12, 2, 20], [9, 18, 7, 22], [9, 31, 11, 29], [9, 27, 5, 13],
			[9, 16, 0, 25], [10, 15, 3, 21], [10, 19, 6, 23],
			[10, 28, 8, 30], [10, 24, 4, 14], [10, 17, 1, 26],
			[11, 14, 0, 23], [11, 16, 4, 21], [11, 25, 9, 27],
			[11, 29, 6, 15], [11, 18, 2, 31]]
	},
	Polyhedron{
		name:      'TruncatedGreatIcosahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: -0.5
			z: 0.927051
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -0.927051
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 0.927051
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -0.927051
		}, Vertex{
			x: -0.5
			y: 0.927051
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.927051
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -0.927051
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -0.927051
			z: 0.0
		}, Vertex{
			x: 0.927051
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.927051
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -0.927051
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -0.927051
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: -1.0
			z: 0.1180340
		}, Vertex{
			x: 0.309017
			y: -1.0
			z: -0.1180340
		}, Vertex{
			x: -0.309017
			y: -1.0
			z: 0.1180340
		}, Vertex{
			x: -0.309017
			y: -1.0
			z: -0.1180340
		}, Vertex{
			x: 0.309017
			y: 1.0
			z: 0.1180340
		}, Vertex{
			x: 0.309017
			y: 1.0
			z: -0.1180340
		}, Vertex{
			x: -0.309017
			y: 1.0
			z: 0.1180340
		}, Vertex{
			x: -0.309017
			y: 1.0
			z: -0.1180340
		}, Vertex{
			x: -1.0
			y: 0.1180340
			z: 0.309017
		}, Vertex{
			x: -1.0
			y: 0.1180340
			z: -0.309017
		}, Vertex{
			x: 1.0
			y: 0.1180340
			z: 0.309017
		}, Vertex{
			x: 1.0
			y: 0.1180340
			z: -0.309017
		}, Vertex{
			x: -1.0
			y: -0.1180340
			z: 0.309017
		}, Vertex{
			x: -1.0
			y: -0.1180340
			z: -0.309017
		}, Vertex{
			x: 1.0
			y: -0.1180340
			z: 0.309017
		}, Vertex{
			x: 1.0
			y: -0.1180340
			z: -0.309017
		}, Vertex{
			x: 0.1180340
			y: 0.309017
			z: -1.0
		}, Vertex{
			x: 0.1180340
			y: 0.309017
			z: 1.0
		}, Vertex{
			x: -0.1180340
			y: 0.309017
			z: -1.0
		}, Vertex{
			x: -0.1180340
			y: 0.309017
			z: 1.0
		}, Vertex{
			x: 0.1180340
			y: -0.309017
			z: -1.0
		}, Vertex{
			x: 0.1180340
			y: -0.309017
			z: 1.0
		}, Vertex{
			x: -0.1180340
			y: -0.309017
			z: -1.0
		}, Vertex{
			x: -0.1180340
			y: -0.309017
			z: 1.0
		}, Vertex{
			x: 0.618034
			y: -0.5
			z: -0.690983
		}, Vertex{
			x: 0.618034
			y: -0.5
			z: 0.690983
		}, Vertex{
			x: -0.618034
			y: -0.5
			z: -0.690983
		}, Vertex{
			x: -0.618034
			y: -0.5
			z: 0.690983
		}, Vertex{
			x: 0.618034
			y: 0.5
			z: -0.690983
		}, Vertex{
			x: 0.618034
			y: 0.5
			z: 0.690983
		}, Vertex{
			x: -0.618034
			y: 0.5
			z: -0.690983
		}, Vertex{
			x: -0.618034
			y: 0.5
			z: 0.690983
		}, Vertex{
			x: -0.5
			y: -0.690983
			z: 0.618034
		}, Vertex{
			x: -0.5
			y: -0.690983
			z: -0.618034
		}, Vertex{
			x: 0.5
			y: -0.690983
			z: 0.618034
		}, Vertex{
			x: 0.5
			y: -0.690983
			z: -0.618034
		}, Vertex{
			x: -0.5
			y: 0.690983
			z: 0.618034
		}, Vertex{
			x: -0.5
			y: 0.690983
			z: -0.618034
		}, Vertex{
			x: 0.5
			y: 0.690983
			z: 0.618034
		}, Vertex{
			x: 0.5
			y: 0.690983
			z: -0.618034
		}, Vertex{
			x: -0.690983
			y: 0.618034
			z: -0.5
		}, Vertex{
			x: -0.690983
			y: 0.618034
			z: 0.5
		}, Vertex{
			x: 0.690983
			y: 0.618034
			z: -0.5
		}, Vertex{
			x: 0.690983
			y: 0.618034
			z: 0.5
		}, Vertex{
			x: -0.690983
			y: -0.618034
			z: -0.5
		}, Vertex{
			x: -0.690983
			y: -0.618034
			z: 0.5
		}, Vertex{
			x: 0.690983
			y: -0.618034
			z: -0.5
		}, Vertex{
			x: 0.690983
			y: -0.618034
			z: 0.5
		}]
		faces:     [[0, 2, 18, 42, 38, 14], [1, 3, 17, 41, 37, 13],
			[2, 0, 12, 36, 40, 16], [3, 1, 15, 39, 43, 19], [4, 5, 23, 47, 45, 21],
			[5, 4, 20, 44, 46, 22], [6, 7, 26, 50, 48, 24], [7, 6, 25, 49, 51, 27],
			[8, 9, 33, 57, 56, 32], [9, 8, 28, 52, 53, 29], [10, 11, 31, 55, 54, 30],
			[11, 10, 34, 58, 59, 35], [12, 44, 20, 52, 28, 36],
			[13, 37, 29, 53, 21, 45], [14, 38, 30, 54, 22, 46],
			[15, 47, 23, 55, 31, 39], [16, 40, 32, 56, 24, 48],
			[17, 49, 25, 57, 33, 41], [18, 50, 26, 58, 34, 42],
			[19, 43, 35, 59, 27, 51], [0, 14, 46, 44, 12], [1, 13, 45, 47, 15],
			[2, 16, 48, 50, 18], [3, 19, 51, 49, 17], [4, 21, 53, 52, 20],
			[5, 22, 54, 55, 23], [6, 24, 56, 57, 25], [7, 27, 59, 58, 26],
			[8, 32, 40, 36, 28], [9, 29, 37, 41, 33], [10, 30, 38, 42, 34],
			[11, 35, 43, 39, 31]]
	},
	Polyhedron{
		name:      'SmallDodecacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: 2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: 0.7834576
			z: 2.051119
		}, Vertex{
			x: 0.0
			y: 0.7834576
			z: -2.051119
		}, Vertex{
			x: 0.0
			y: -0.7834576
			z: 2.051119
		}, Vertex{
			x: 0.0
			y: -0.7834576
			z: -2.051119
		}, Vertex{
			x: 2.051119
			y: 0.0
			z: 0.7834576
		}, Vertex{
			x: 2.051119
			y: 0.0
			z: -0.7834576
		}, Vertex{
			x: -2.051119
			y: 0.0
			z: 0.7834576
		}, Vertex{
			x: -2.051119
			y: 0.0
			z: -0.7834576
		}, Vertex{
			x: 0.7834576
			y: 2.051119
			z: 0.0
		}, Vertex{
			x: 0.7834576
			y: -2.051119
			z: 0.0
		}, Vertex{
			x: -0.7834576
			y: 2.051119
			z: 0.0
		}, Vertex{
			x: -0.7834576
			y: -2.051119
			z: 0.0
		}, Vertex{
			x: 1.206011
			y: 0.0
			z: 1.951367
		}, Vertex{
			x: 1.206011
			y: 0.0
			z: -1.951367
		}, Vertex{
			x: -1.206011
			y: 0.0
			z: 1.951367
		}, Vertex{
			x: -1.206011
			y: 0.0
			z: -1.951367
		}, Vertex{
			x: 1.951367
			y: 1.206011
			z: 0.0
		}, Vertex{
			x: 1.951367
			y: -1.206011
			z: 0.0
		}, Vertex{
			x: -1.951367
			y: 1.206011
			z: 0.0
		}, Vertex{
			x: -1.951367
			y: -1.206011
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.951367
			z: 1.206011
		}, Vertex{
			x: 0.0
			y: 1.951367
			z: -1.206011
		}, Vertex{
			x: 0.0
			y: -1.951367
			z: 1.206011
		}, Vertex{
			x: 0.0
			y: -1.951367
			z: -1.206011
		}, Vertex{
			x: 1.267661
			y: 1.267661
			z: 1.267661
		}, Vertex{
			x: 1.267661
			y: 1.267661
			z: -1.267661
		}, Vertex{
			x: 1.267661
			y: -1.267661
			z: 1.267661
		}, Vertex{
			x: 1.267661
			y: -1.267661
			z: -1.267661
		}, Vertex{
			x: -1.267661
			y: 1.267661
			z: 1.267661
		}, Vertex{
			x: -1.267661
			y: 1.267661
			z: -1.267661
		}, Vertex{
			x: -1.267661
			y: -1.267661
			z: 1.267661
		}, Vertex{
			x: -1.267661
			y: -1.267661
			z: -1.267661
		}]
		faces:     [[24, 2, 14, 10], [24, 10, 38, 5], [24, 5, 16, 4],
			[24, 4, 36, 8], [24, 8, 12, 2], [25, 3, 13, 9], [25, 9, 37, 4],
			[25, 4, 17, 5], [25, 5, 39, 11], [25, 11, 15, 3],
			[26, 0, 12, 8], [26, 8, 40, 6], [26, 6, 18, 7], [26, 7, 42, 10],
			[26, 10, 14, 0], [27, 1, 15, 11], [27, 11, 43, 7],
			[27, 7, 19, 6], [27, 6, 41, 9], [27, 9, 13, 1], [28, 0, 16, 5],
			[28, 5, 17, 1], [28, 1, 37, 9], [28, 9, 20, 8], [28, 8, 36, 0],
			[29, 0, 38, 10], [29, 10, 21, 11], [29, 11, 39, 1],
			[29, 1, 17, 4], [29, 4, 16, 0], [30, 2, 40, 8], [30, 8, 22, 9],
			[30, 9, 41, 3], [30, 3, 19, 7], [30, 7, 18, 2], [31, 2, 18, 6],
			[31, 6, 19, 3], [31, 3, 43, 11], [31, 11, 23, 10],
			[31, 10, 42, 2], [32, 0, 36, 4], [32, 4, 20, 9], [32, 9, 22, 6],
			[32, 6, 40, 2], [32, 2, 12, 0], [33, 1, 13, 3], [33, 3, 41, 6],
			[33, 6, 22, 8], [33, 8, 20, 4], [33, 4, 37, 1], [34, 0, 14, 2],
			[34, 2, 42, 7], [34, 7, 23, 11], [34, 11, 21, 5],
			[34, 5, 38, 0], [35, 1, 39, 5], [35, 5, 21, 10], [35, 10, 23, 7],
			[35, 7, 43, 3], [35, 3, 15, 1]]
	},
	Polyhedron{
		name:      'GreatDitrigonalDodecicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.809017
			y: -0.5
			z: 0.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: -0.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: 0.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: -0.618034
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: 0.618034
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: -0.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: 0.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: -0.618034
		}, Vertex{
			x: -0.5
			y: 0.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: 0.618034
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: 0.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: 0.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: -0.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: -0.618034
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: -0.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: -0.618034
			z: -0.809017
		}, Vertex{
			x: 0.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: 0.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: -0.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: 0.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: 0.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: -0.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: 1.118034
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: -1.118034
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: -1.118034
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: 1.118034
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: -1.118034
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: 1.118034
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: -1.118034
		}, Vertex{
			x: -0.1909830
			y: 1.118034
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: 1.118034
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: -1.118034
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: -1.118034
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -1.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: -1.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: -1.0
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: -1.0
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: 1.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: 1.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: 1.0
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: 1.0
			z: 0.1909830
		}, Vertex{
			x: -1.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: -1.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: 1.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: 1.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: -1.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: -1.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: 1.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: 1.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: -1.0
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: 1.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: -1.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: 1.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: -1.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: 1.0
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: -1.0
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: 1.0
		}]
		faces:     [[0, 4, 30, 14, 51, 59, 55, 47, 10, 28], [0, 38, 46, 47, 39, 1, 25, 21, 20, 24],
			[2, 26, 22, 23, 27, 3, 37, 45, 44, 36], [2, 28, 8, 45, 53, 57, 49, 12, 30, 6],
			[5, 1, 29, 11, 46, 54, 58, 50, 15, 31], [5, 43, 51, 50, 42, 4, 24, 16, 17, 25],
			[7, 27, 19, 18, 26, 6, 40, 48, 49, 41], [7, 31, 13, 48, 56, 52, 44, 9, 29, 3],
			[33, 11, 9, 32, 16, 56, 40, 42, 58, 18], [33, 19, 59, 43, 41, 57, 17, 32, 8, 10],
			[34, 13, 15, 35, 22, 54, 38, 36, 52, 20], [34, 21, 53, 37, 39, 55, 23, 35, 14, 12],
			[24, 20, 52, 56, 16], [25, 17, 57, 53, 21], [26, 18, 58, 54, 22],
			[27, 23, 55, 59, 19], [28, 2, 36, 38, 0], [29, 1, 39, 37, 3],
			[30, 4, 42, 40, 6], [31, 7, 41, 43, 5], [32, 9, 44, 45, 8],
			[33, 10, 47, 46, 11], [34, 12, 49, 48, 13], [35, 15, 50, 51, 14],
			[24, 4, 0], [25, 1, 5], [26, 2, 6], [27, 7, 3], [28, 10, 8],
			[29, 9, 11], [30, 12, 14], [31, 15, 13], [32, 17, 16],
			[33, 18, 19], [34, 20, 21], [35, 23, 22], [36, 44, 52],
			[37, 53, 45], [38, 54, 46], [39, 47, 55], [40, 56, 48],
			[41, 49, 57], [42, 50, 58], [43, 59, 51]]
	},
	Polyhedron{
		name:      'GreatDisdyakisTriacontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: -1.075711
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.075711
		}, Vertex{
			x: 0.0
			y: -1.075711
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.075711
			z: 0.0
		}, Vertex{
			x: -1.075711
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 1.075711
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 3.618034
			y: 0.0
			z: 1.381966
		}, Vertex{
			x: 3.618034
			y: 0.0
			z: -1.381966
		}, Vertex{
			x: -3.618034
			y: 0.0
			z: 1.381966
		}, Vertex{
			x: -3.618034
			y: 0.0
			z: -1.381966
		}, Vertex{
			x: 0.0
			y: 1.381966
			z: 3.618034
		}, Vertex{
			x: 0.0
			y: 1.381966
			z: -3.618034
		}, Vertex{
			x: 0.0
			y: -1.381966
			z: 3.618034
		}, Vertex{
			x: 0.0
			y: -1.381966
			z: -3.618034
		}, Vertex{
			x: 1.381966
			y: 3.618034
			z: 0.0
		}, Vertex{
			x: -1.381966
			y: 3.618034
			z: 0.0
		}, Vertex{
			x: 1.381966
			y: -3.618034
			z: 0.0
		}, Vertex{
			x: -1.381966
			y: -3.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.8291796
			z: -0.5124612
		}, Vertex{
			x: 0.0
			y: 0.8291796
			z: 0.5124612
		}, Vertex{
			x: 0.0
			y: -0.8291796
			z: -0.5124612
		}, Vertex{
			x: 0.0
			y: -0.8291796
			z: 0.5124612
		}, Vertex{
			x: 0.8291796
			y: -0.5124612
			z: 0.0
		}, Vertex{
			x: -0.8291796
			y: -0.5124612
			z: 0.0
		}, Vertex{
			x: 0.8291796
			y: 0.5124612
			z: 0.0
		}, Vertex{
			x: -0.8291796
			y: 0.5124612
			z: 0.0
		}, Vertex{
			x: -0.5124612
			y: 0.0
			z: 0.8291796
		}, Vertex{
			x: -0.5124612
			y: 0.0
			z: -0.8291796
		}, Vertex{
			x: 0.5124612
			y: 0.0
			z: 0.8291796
		}, Vertex{
			x: 0.5124612
			y: 0.0
			z: -0.8291796
		}, Vertex{
			x: -0.5378553
			y: 0.8702681
			z: 0.3324128
		}, Vertex{
			x: -0.5378553
			y: 0.8702681
			z: -0.3324128
		}, Vertex{
			x: 0.5378553
			y: 0.8702681
			z: 0.3324128
		}, Vertex{
			x: 0.5378553
			y: 0.8702681
			z: -0.3324128
		}, Vertex{
			x: -0.5378553
			y: -0.8702681
			z: 0.3324128
		}, Vertex{
			x: -0.5378553
			y: -0.8702681
			z: -0.3324128
		}, Vertex{
			x: 0.5378553
			y: -0.8702681
			z: 0.3324128
		}, Vertex{
			x: 0.5378553
			y: -0.8702681
			z: -0.3324128
		}, Vertex{
			x: 0.8702681
			y: 0.3324128
			z: -0.5378553
		}, Vertex{
			x: 0.8702681
			y: 0.3324128
			z: 0.5378553
		}, Vertex{
			x: -0.8702681
			y: 0.3324128
			z: -0.5378553
		}, Vertex{
			x: -0.8702681
			y: 0.3324128
			z: 0.5378553
		}, Vertex{
			x: 0.8702681
			y: -0.3324128
			z: -0.5378553
		}, Vertex{
			x: 0.8702681
			y: -0.3324128
			z: 0.5378553
		}, Vertex{
			x: -0.8702681
			y: -0.3324128
			z: -0.5378553
		}, Vertex{
			x: -0.8702681
			y: -0.3324128
			z: 0.5378553
		}, Vertex{
			x: 0.3324128
			y: -0.5378553
			z: 0.8702681
		}, Vertex{
			x: 0.3324128
			y: -0.5378553
			z: -0.8702681
		}, Vertex{
			x: -0.3324128
			y: -0.5378553
			z: 0.8702681
		}, Vertex{
			x: -0.3324128
			y: -0.5378553
			z: -0.8702681
		}, Vertex{
			x: 0.3324128
			y: 0.5378553
			z: 0.8702681
		}, Vertex{
			x: 0.3324128
			y: 0.5378553
			z: -0.8702681
		}, Vertex{
			x: -0.3324128
			y: 0.5378553
			z: 0.8702681
		}, Vertex{
			x: -0.3324128
			y: 0.5378553
			z: -0.8702681
		}, Vertex{
			x: -2.236068
			y: -2.236068
			z: -2.236068
		}, Vertex{
			x: -2.236068
			y: -2.236068
			z: 2.236068
		}, Vertex{
			x: 2.236068
			y: -2.236068
			z: -2.236068
		}, Vertex{
			x: 2.236068
			y: -2.236068
			z: 2.236068
		}, Vertex{
			x: -2.236068
			y: 2.236068
			z: -2.236068
		}, Vertex{
			x: -2.236068
			y: 2.236068
			z: 2.236068
		}, Vertex{
			x: 2.236068
			y: 2.236068
			z: -2.236068
		}, Vertex{
			x: 2.236068
			y: 2.236068
			z: 2.236068
		}]
		faces:     [[18, 0, 8], [18, 8, 32], [18, 32, 56], [18, 56, 40],
			[18, 40, 10], [18, 10, 38], [18, 38, 54], [18, 54, 30],
			[18, 30, 6], [18, 6, 0], [19, 1, 7], [19, 7, 31],
			[19, 31, 55], [19, 55, 39], [19, 39, 11], [19, 11, 41],
			[19, 41, 57], [19, 57, 33], [19, 33, 9], [19, 9, 1],
			[20, 0, 6], [20, 6, 34], [20, 34, 58], [20, 58, 42],
			[20, 42, 12], [20, 12, 44], [20, 44, 60], [20, 60, 36],
			[20, 36, 8], [20, 8, 0], [21, 1, 9], [21, 9, 37],
			[21, 37, 61], [21, 61, 45], [21, 45, 13], [21, 13, 43],
			[21, 43, 59], [21, 59, 35], [21, 35, 7], [21, 7, 1],
			[22, 2, 11], [22, 11, 39], [22, 39, 55], [22, 55, 47],
			[22, 47, 14], [22, 14, 46], [22, 46, 54], [22, 54, 38],
			[22, 38, 10], [22, 10, 2], [23, 2, 10], [23, 10, 40],
			[23, 40, 56], [23, 56, 48], [23, 48, 15], [23, 15, 49],
			[23, 49, 57], [23, 57, 41], [23, 41, 11], [23, 11, 2],
			[24, 3, 12], [24, 12, 42], [24, 42, 58], [24, 58, 50],
			[24, 50, 16], [24, 16, 51], [24, 51, 59], [24, 59, 43],
			[24, 43, 13], [24, 13, 3], [25, 3, 13], [25, 13, 45],
			[25, 45, 61], [25, 61, 53], [25, 53, 17], [25, 17, 52],
			[25, 52, 60], [25, 60, 44], [25, 44, 12], [25, 12, 3],
			[26, 4, 16], [26, 16, 50], [26, 50, 58], [26, 58, 34],
			[26, 34, 6], [26, 6, 30], [26, 30, 54], [26, 54, 46],
			[26, 46, 14], [26, 14, 4], [27, 4, 14], [27, 14, 47],
			[27, 47, 55], [27, 55, 31], [27, 31, 7], [27, 7, 35],
			[27, 35, 59], [27, 59, 51], [27, 51, 16], [27, 16, 4],
			[28, 5, 15], [28, 15, 48], [28, 48, 56], [28, 56, 32],
			[28, 32, 8], [28, 8, 36], [28, 36, 60], [28, 60, 52],
			[28, 52, 17], [28, 17, 5], [29, 5, 17], [29, 17, 53],
			[29, 53, 61], [29, 61, 37], [29, 37, 9], [29, 9, 33],
			[29, 33, 57], [29, 57, 49], [29, 49, 15], [29, 15, 5]]
	},
	Polyhedron{
		name:      'GreatHexacronicIcositetrahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: -0.5857865
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 0.5857865
		}, Vertex{
			x: -0.5857865
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.5857865
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.5857865
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.5857865
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.414214
			z: 0.0
		}, Vertex{
			x: -0.3693981
			y: -0.3693981
			z: -0.3693981
		}, Vertex{
			x: -0.3693981
			y: -0.3693981
			z: 0.3693981
		}, Vertex{
			x: -0.3693981
			y: 0.3693981
			z: -0.3693981
		}, Vertex{
			x: -0.3693981
			y: 0.3693981
			z: 0.3693981
		}, Vertex{
			x: 0.3693981
			y: -0.3693981
			z: -0.3693981
		}, Vertex{
			x: 0.3693981
			y: -0.3693981
			z: 0.3693981
		}, Vertex{
			x: 0.3693981
			y: 0.3693981
			z: -0.3693981
		}, Vertex{
			x: 0.3693981
			y: 0.3693981
			z: 0.3693981
		}]
		faces:     [[12, 0, 8, 4], [12, 4, 6, 2], [12, 2, 10, 0],
			[13, 1, 10, 2], [13, 2, 7, 4], [13, 4, 8, 1], [14, 0, 11, 2],
			[14, 2, 6, 5], [14, 5, 8, 0], [15, 1, 8, 5], [15, 5, 7, 2],
			[15, 2, 11, 1], [16, 0, 10, 3], [16, 3, 6, 4], [16, 4, 9, 0],
			[17, 1, 9, 4], [17, 4, 7, 3], [17, 3, 10, 1], [18, 0, 9, 5],
			[18, 5, 6, 3], [18, 3, 11, 0], [19, 1, 11, 3], [19, 3, 7, 5],
			[19, 5, 9, 1]]
	},
	Polyhedron{
		name:      'GreatRhombidodecacron'
		vertexes_: [Vertex{
			x: 0.0
			y: -0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: -0.3819660
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: -0.3819660
		}, Vertex{
			x: -0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -2.236068
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 2.236068
		}, Vertex{
			x: 0.0
			y: -2.236068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.236068
			z: 0.0
		}, Vertex{
			x: -2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: -1.809017
		}]
		faces:     [[0, 14, 5, 26], [0, 36, 10, 28], [0, 24, 2, 20],
			[0, 22, 8, 12], [0, 34, 4, 18], [1, 14, 4, 29], [1, 37, 5, 21],
			[1, 25, 11, 13], [1, 23, 3, 19], [1, 35, 9, 27], [2, 15, 6, 32],
			[2, 38, 8, 30], [2, 18, 0, 22], [2, 20, 10, 12], [2, 40, 7, 24],
			[3, 15, 7, 31], [3, 39, 6, 23], [3, 19, 9, 13], [3, 21, 1, 25],
			[3, 41, 11, 33], [4, 16, 9, 34], [4, 19, 1, 35], [4, 29, 5, 27],
			[4, 28, 0, 14], [4, 18, 8, 26], [5, 17, 10, 37], [5, 20, 0, 36],
			[5, 26, 4, 28], [5, 27, 1, 14], [5, 21, 11, 29], [6, 16, 8, 39],
			[6, 22, 2, 38], [6, 32, 7, 30], [6, 33, 3, 15], [6, 23, 9, 31],
			[7, 17, 11, 40], [7, 25, 3, 41], [7, 31, 6, 33], [7, 30, 2, 15],
			[7, 24, 10, 32], [8, 12, 2, 18], [8, 30, 6, 22], [8, 39, 9, 38],
			[8, 35, 4, 16], [8, 26, 0, 34], [9, 13, 1, 23], [9, 27, 4, 19],
			[9, 34, 8, 35], [9, 38, 6, 16], [9, 31, 3, 39], [10, 12, 0, 24],
			[10, 28, 5, 20], [10, 37, 11, 36], [10, 41, 7, 17],
			[10, 32, 2, 40], [11, 13, 3, 21], [11, 33, 7, 25],
			[11, 40, 10, 41], [11, 36, 5, 17], [11, 29, 1, 37]]
	},
	Polyhedron{
		name:      'TriakisIcosahedron'
		vertexes_: [Vertex{
			x: 1.809017
			y: 0.0
			z: 2.927051
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -2.927051
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 2.927051
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -2.927051
		}, Vertex{
			x: 2.927051
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 2.927051
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -2.927051
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -2.927051
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.927051
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 2.927051
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -2.927051
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -2.927051
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: 1.049553
			z: 2.747766
		}, Vertex{
			x: 0.0
			y: 1.049553
			z: -2.747766
		}, Vertex{
			x: 0.0
			y: -1.049553
			z: 2.747766
		}, Vertex{
			x: 0.0
			y: -1.049553
			z: -2.747766
		}, Vertex{
			x: 2.747766
			y: 0.0
			z: 1.049553
		}, Vertex{
			x: 2.747766
			y: 0.0
			z: -1.049553
		}, Vertex{
			x: -2.747766
			y: 0.0
			z: 1.049553
		}, Vertex{
			x: -2.747766
			y: 0.0
			z: -1.049553
		}, Vertex{
			x: 1.049553
			y: 2.747766
			z: 0.0
		}, Vertex{
			x: 1.049553
			y: -2.747766
			z: 0.0
		}, Vertex{
			x: -1.049553
			y: 2.747766
			z: 0.0
		}, Vertex{
			x: -1.049553
			y: -2.747766
			z: 0.0
		}, Vertex{
			x: 1.698213
			y: 1.698213
			z: 1.698213
		}, Vertex{
			x: 1.698213
			y: 1.698213
			z: -1.698213
		}, Vertex{
			x: 1.698213
			y: -1.698213
			z: 1.698213
		}, Vertex{
			x: 1.698213
			y: -1.698213
			z: -1.698213
		}, Vertex{
			x: -1.698213
			y: 1.698213
			z: 1.698213
		}, Vertex{
			x: -1.698213
			y: 1.698213
			z: -1.698213
		}, Vertex{
			x: -1.698213
			y: -1.698213
			z: 1.698213
		}, Vertex{
			x: -1.698213
			y: -1.698213
			z: -1.698213
		}]
		faces:     [[12, 0, 8], [12, 8, 2], [12, 2, 0], [13, 1, 3],
			[13, 3, 9], [13, 9, 1], [14, 0, 2], [14, 2, 10], [14, 10, 0],
			[15, 1, 11], [15, 11, 3], [15, 3, 1], [16, 0, 5],
			[16, 5, 4], [16, 4, 0], [17, 1, 4], [17, 4, 5], [17, 5, 1],
			[18, 2, 6], [18, 6, 7], [18, 7, 2], [19, 3, 7], [19, 7, 6],
			[19, 6, 3], [20, 4, 9], [20, 9, 8], [20, 8, 4], [21, 5, 10],
			[21, 10, 11], [21, 11, 5], [22, 6, 8], [22, 8, 9],
			[22, 9, 6], [23, 7, 11], [23, 11, 10], [23, 10, 7],
			[24, 0, 4], [24, 4, 8], [24, 8, 0], [25, 1, 9], [25, 9, 4],
			[25, 4, 1], [26, 0, 10], [26, 10, 5], [26, 5, 0],
			[27, 1, 5], [27, 5, 11], [27, 11, 1], [28, 2, 8],
			[28, 8, 6], [28, 6, 2], [29, 3, 6], [29, 6, 9], [29, 9, 3],
			[30, 2, 7], [30, 7, 10], [30, 10, 2], [31, 3, 11],
			[31, 11, 7], [31, 7, 3]]
	},
	Polyhedron{
		name:      'GreatRhombihexahedron'
		vertexes_: [Vertex{
			x: -0.5
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: 0.5
		}]
		faces:     [[0, 2, 18, 19, 3, 1, 17, 16], [0, 8, 9, 1, 5, 13, 12, 4],
			[14, 15, 7, 3, 11, 10, 2, 6], [14, 22, 18, 10, 8, 16, 20, 12],
			[21, 5, 7, 23, 22, 6, 4, 20], [21, 17, 9, 11, 19, 23, 15, 13],
			[0, 2, 10, 8], [0, 16, 20, 4], [7, 3, 19, 23], [7, 15, 13, 5],
			[11, 3, 1, 9], [11, 10, 18, 19], [12, 14, 6, 4], [12, 20, 21, 13],
			[17, 1, 5, 21], [17, 16, 8, 9], [22, 14, 15, 23],
			[22, 18, 2, 6]]
	},
	Polyhedron{
		name:      'TruncatedGreatDodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.0
			z: 1.809017
		}, Vertex{
			x: 0.5
			y: 0.0
			z: -1.809017
		}, Vertex{
			x: -0.5
			y: 0.0
			z: 1.809017
		}, Vertex{
			x: -0.5
			y: 0.0
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.5
			z: 0.0
		}, Vertex{
			x: 1.809017
			y: -0.5
			z: 0.0
		}, Vertex{
			x: -1.809017
			y: 0.5
			z: 0.0
		}, Vertex{
			x: -1.809017
			y: -0.5
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.809017
			z: 0.5
		}, Vertex{
			x: 0.0
			y: 1.809017
			z: -0.5
		}, Vertex{
			x: 0.0
			y: -1.809017
			z: 0.5
		}, Vertex{
			x: 0.0
			y: -1.809017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: 1.618034
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: -1.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: 1.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: -1.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: 1.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: -1.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: 1.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: 1.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: 1.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: 1.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: -1.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: -1.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: -1.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: -1.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: 1.618034
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: -1.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: -1.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: 1.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: 1.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: -1.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: -1.618034
			z: -0.809017
		}, Vertex{
			x: 1.309017
			y: 0.309017
			z: 1.309017
		}, Vertex{
			x: 1.309017
			y: 0.309017
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: -0.309017
			z: 1.309017
		}, Vertex{
			x: 1.309017
			y: -0.309017
			z: -1.309017
		}, Vertex{
			x: -1.309017
			y: 0.309017
			z: 1.309017
		}, Vertex{
			x: -1.309017
			y: 0.309017
			z: -1.309017
		}, Vertex{
			x: -1.309017
			y: -0.309017
			z: 1.309017
		}, Vertex{
			x: -1.309017
			y: -0.309017
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.309017
			z: 0.309017
		}, Vertex{
			x: 1.309017
			y: 1.309017
			z: -0.309017
		}, Vertex{
			x: 1.309017
			y: -1.309017
			z: 0.309017
		}, Vertex{
			x: 1.309017
			y: -1.309017
			z: -0.309017
		}, Vertex{
			x: -1.309017
			y: 1.309017
			z: 0.309017
		}, Vertex{
			x: -1.309017
			y: 1.309017
			z: -0.309017
		}, Vertex{
			x: -1.309017
			y: -1.309017
			z: 0.309017
		}, Vertex{
			x: -1.309017
			y: -1.309017
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: 1.309017
			z: 1.309017
		}, Vertex{
			x: 0.309017
			y: 1.309017
			z: -1.309017
		}, Vertex{
			x: 0.309017
			y: -1.309017
			z: 1.309017
		}, Vertex{
			x: 0.309017
			y: -1.309017
			z: -1.309017
		}, Vertex{
			x: -0.309017
			y: 1.309017
			z: 1.309017
		}, Vertex{
			x: -0.309017
			y: 1.309017
			z: -1.309017
		}, Vertex{
			x: -0.309017
			y: -1.309017
			z: 1.309017
		}, Vertex{
			x: -0.309017
			y: -1.309017
			z: -1.309017
		}]
		faces:     [[0, 2, 42, 26, 51, 35, 31, 47, 22, 38], [1, 3, 41, 25, 48, 32, 28, 44, 21, 37],
			[2, 0, 36, 20, 45, 29, 33, 49, 24, 40], [3, 1, 39, 23, 46, 30, 34, 50, 27, 43],
			[4, 5, 47, 31, 59, 19, 17, 57, 29, 45], [5, 4, 44, 28, 56, 16, 18, 58, 30, 46],
			[6, 7, 50, 34, 54, 14, 12, 52, 32, 48], [7, 6, 49, 33, 53, 13, 15, 55, 35, 51],
			[8, 9, 57, 17, 43, 27, 26, 42, 16, 56], [9, 8, 52, 12, 38, 22, 23, 39, 13, 53],
			[10, 11, 55, 15, 37, 21, 20, 36, 14, 54], [11, 10, 58, 18, 40, 24, 25, 41, 19, 59],
			[0, 38, 12, 14, 36], [1, 37, 15, 13, 39], [2, 40, 18, 16, 42],
			[3, 43, 17, 19, 41], [4, 45, 20, 21, 44], [5, 46, 23, 22, 47],
			[6, 48, 25, 24, 49], [7, 51, 26, 27, 50], [8, 56, 28, 32, 52],
			[9, 53, 33, 29, 57], [10, 54, 34, 30, 58], [11, 59, 31, 35, 55]]
	},
	Polyhedron{
		name:      'TruncatedIcosidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 3.736068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -3.736068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 3.736068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -3.736068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 3.736068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -3.736068
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 3.736068
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -3.736068
		}, Vertex{
			x: 3.736068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 3.736068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 3.736068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 3.736068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -3.736068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -3.736068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -3.736068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -3.736068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 3.736068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 3.736068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -3.736068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -3.736068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 3.736068
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 3.736068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -3.736068
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -3.736068
			z: -0.5
		}, Vertex{
			x: 1.0
			y: 1.309017
			z: 3.427051
		}, Vertex{
			x: 1.0
			y: 1.309017
			z: -3.427051
		}, Vertex{
			x: 1.0
			y: -1.309017
			z: 3.427051
		}, Vertex{
			x: 1.0
			y: -1.309017
			z: -3.427051
		}, Vertex{
			x: -1.0
			y: 1.309017
			z: 3.427051
		}, Vertex{
			x: -1.0
			y: 1.309017
			z: -3.427051
		}, Vertex{
			x: -1.0
			y: -1.309017
			z: 3.427051
		}, Vertex{
			x: -1.0
			y: -1.309017
			z: -3.427051
		}, Vertex{
			x: 3.427051
			y: 1.0
			z: 1.309017
		}, Vertex{
			x: 3.427051
			y: 1.0
			z: -1.309017
		}, Vertex{
			x: 3.427051
			y: -1.0
			z: 1.309017
		}, Vertex{
			x: 3.427051
			y: -1.0
			z: -1.309017
		}, Vertex{
			x: -3.427051
			y: 1.0
			z: 1.309017
		}, Vertex{
			x: -3.427051
			y: 1.0
			z: -1.309017
		}, Vertex{
			x: -3.427051
			y: -1.0
			z: 1.309017
		}, Vertex{
			x: -3.427051
			y: -1.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 3.427051
			z: 1.0
		}, Vertex{
			x: 1.309017
			y: 3.427051
			z: -1.0
		}, Vertex{
			x: 1.309017
			y: -3.427051
			z: 1.0
		}, Vertex{
			x: 1.309017
			y: -3.427051
			z: -1.0
		}, Vertex{
			x: -1.309017
			y: 3.427051
			z: 1.0
		}, Vertex{
			x: -1.309017
			y: 3.427051
			z: -1.0
		}, Vertex{
			x: -1.309017
			y: -3.427051
			z: 1.0
		}, Vertex{
			x: -1.309017
			y: -3.427051
			z: -1.0
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: 3.118034
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: -3.118034
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: 3.118034
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: -3.118034
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: 3.118034
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: -3.118034
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: 3.118034
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: -3.118034
		}, Vertex{
			x: 3.118034
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: 3.118034
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: 3.118034
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: 3.118034
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: -3.118034
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: -3.118034
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: -3.118034
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: -3.118034
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: 2.118034
			y: 3.118034
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: 3.118034
			z: -0.5
		}, Vertex{
			x: 2.118034
			y: -3.118034
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: -3.118034
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: 3.118034
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: 3.118034
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: -3.118034
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: -3.118034
			z: -0.5
		}, Vertex{
			x: 1.809017
			y: 1.618034
			z: 2.927051
		}, Vertex{
			x: 1.809017
			y: 1.618034
			z: -2.927051
		}, Vertex{
			x: 1.809017
			y: -1.618034
			z: 2.927051
		}, Vertex{
			x: 1.809017
			y: -1.618034
			z: -2.927051
		}, Vertex{
			x: -1.809017
			y: 1.618034
			z: 2.927051
		}, Vertex{
			x: -1.809017
			y: 1.618034
			z: -2.927051
		}, Vertex{
			x: -1.809017
			y: -1.618034
			z: 2.927051
		}, Vertex{
			x: -1.809017
			y: -1.618034
			z: -2.927051
		}, Vertex{
			x: 2.927051
			y: 1.809017
			z: 1.618034
		}, Vertex{
			x: 2.927051
			y: 1.809017
			z: -1.618034
		}, Vertex{
			x: 2.927051
			y: -1.809017
			z: 1.618034
		}, Vertex{
			x: 2.927051
			y: -1.809017
			z: -1.618034
		}, Vertex{
			x: -2.927051
			y: 1.809017
			z: 1.618034
		}, Vertex{
			x: -2.927051
			y: 1.809017
			z: -1.618034
		}, Vertex{
			x: -2.927051
			y: -1.809017
			z: 1.618034
		}, Vertex{
			x: -2.927051
			y: -1.809017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 2.927051
			z: 1.809017
		}, Vertex{
			x: 1.618034
			y: 2.927051
			z: -1.809017
		}, Vertex{
			x: 1.618034
			y: -2.927051
			z: 1.809017
		}, Vertex{
			x: 1.618034
			y: -2.927051
			z: -1.809017
		}, Vertex{
			x: -1.618034
			y: 2.927051
			z: 1.809017
		}, Vertex{
			x: -1.618034
			y: 2.927051
			z: -1.809017
		}, Vertex{
			x: -1.618034
			y: -2.927051
			z: 1.809017
		}, Vertex{
			x: -1.618034
			y: -2.927051
			z: -1.809017
		}, Vertex{
			x: 1.309017
			y: 2.427051
			z: 2.618034
		}, Vertex{
			x: 1.309017
			y: 2.427051
			z: -2.618034
		}, Vertex{
			x: 1.309017
			y: -2.427051
			z: 2.618034
		}, Vertex{
			x: 1.309017
			y: -2.427051
			z: -2.618034
		}, Vertex{
			x: -1.309017
			y: 2.427051
			z: 2.618034
		}, Vertex{
			x: -1.309017
			y: 2.427051
			z: -2.618034
		}, Vertex{
			x: -1.309017
			y: -2.427051
			z: 2.618034
		}, Vertex{
			x: -1.309017
			y: -2.427051
			z: -2.618034
		}, Vertex{
			x: 2.618034
			y: 1.309017
			z: 2.427051
		}, Vertex{
			x: 2.618034
			y: 1.309017
			z: -2.427051
		}, Vertex{
			x: 2.618034
			y: -1.309017
			z: 2.427051
		}, Vertex{
			x: 2.618034
			y: -1.309017
			z: -2.427051
		}, Vertex{
			x: -2.618034
			y: 1.309017
			z: 2.427051
		}, Vertex{
			x: -2.618034
			y: 1.309017
			z: -2.427051
		}, Vertex{
			x: -2.618034
			y: -1.309017
			z: 2.427051
		}, Vertex{
			x: -2.618034
			y: -1.309017
			z: -2.427051
		}, Vertex{
			x: 2.427051
			y: 2.618034
			z: 1.309017
		}, Vertex{
			x: 2.427051
			y: 2.618034
			z: -1.309017
		}, Vertex{
			x: 2.427051
			y: -2.618034
			z: 1.309017
		}, Vertex{
			x: 2.427051
			y: -2.618034
			z: -1.309017
		}, Vertex{
			x: -2.427051
			y: 2.618034
			z: 1.309017
		}, Vertex{
			x: -2.427051
			y: 2.618034
			z: -1.309017
		}, Vertex{
			x: -2.427051
			y: -2.618034
			z: 1.309017
		}, Vertex{
			x: -2.427051
			y: -2.618034
			z: -1.309017
		}]
		faces:     [[0, 2, 26, 74, 106, 58, 56, 104, 72, 24],
			[1, 25, 73, 105, 57, 59, 107, 75, 27, 3], [4, 28, 76, 108, 60, 62, 110, 78, 30, 6],
			[5, 7, 31, 79, 111, 63, 61, 109, 77, 29], [8, 9, 33, 81, 113, 65, 64, 112, 80, 32],
			[10, 34, 82, 114, 66, 67, 115, 83, 35, 11], [12, 36, 84, 116, 68, 69, 117, 85, 37, 13],
			[14, 15, 39, 87, 119, 71, 70, 118, 86, 38], [16, 20, 44, 92, 100, 52, 48, 96, 88, 40],
			[17, 41, 89, 97, 49, 53, 101, 93, 45, 21], [18, 42, 90, 98, 50, 54, 102, 94, 46, 22],
			[19, 23, 47, 95, 103, 55, 51, 99, 91, 43], [0, 24, 48, 52, 28, 4],
			[1, 5, 29, 53, 49, 25], [2, 6, 30, 54, 50, 26], [3, 27, 51, 55, 31, 7],
			[8, 32, 56, 58, 34, 10], [9, 11, 35, 59, 57, 33],
			[12, 14, 38, 62, 60, 36], [13, 37, 61, 63, 39, 15],
			[16, 40, 64, 65, 41, 17], [18, 19, 43, 67, 66, 42],
			[20, 21, 45, 69, 68, 44], [22, 46, 70, 71, 47, 23],
			[72, 104, 80, 112, 88, 96], [73, 97, 89, 113, 81, 105],
			[74, 98, 90, 114, 82, 106], [75, 107, 83, 115, 91, 99],
			[76, 100, 92, 116, 84, 108], [77, 109, 85, 117, 93, 101],
			[78, 110, 86, 118, 94, 102], [79, 103, 95, 119, 87, 111],
			[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9], [12, 13, 15, 14],
			[16, 17, 21, 20], [18, 22, 23, 19], [24, 72, 96, 48],
			[25, 49, 97, 73], [26, 50, 98, 74], [27, 75, 99, 51],
			[28, 52, 100, 76], [29, 77, 101, 53], [30, 78, 102, 54],
			[31, 55, 103, 79], [32, 80, 104, 56], [33, 57, 105, 81],
			[34, 58, 106, 82], [35, 83, 107, 59], [36, 60, 108, 84],
			[37, 85, 109, 61], [38, 86, 110, 62], [39, 63, 111, 87],
			[40, 88, 112, 64], [41, 65, 113, 89], [42, 66, 114, 90],
			[43, 91, 115, 67], [44, 68, 116, 92], [45, 93, 117, 69],
			[46, 94, 118, 70], [47, 71, 119, 95]]
	},
	Polyhedron{
		name:      'DisdyakisTriacontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 3.802983
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -3.802983
		}, Vertex{
			x: 3.802983
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -3.802983
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 3.802983
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -3.802983
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.381966
			z: 3.618034
		}, Vertex{
			x: 0.0
			y: 1.381966
			z: -3.618034
		}, Vertex{
			x: 0.0
			y: -1.381966
			z: 3.618034
		}, Vertex{
			x: 0.0
			y: -1.381966
			z: -3.618034
		}, Vertex{
			x: 3.618034
			y: 0.0
			z: 1.381966
		}, Vertex{
			x: 3.618034
			y: 0.0
			z: -1.381966
		}, Vertex{
			x: -3.618034
			y: 0.0
			z: 1.381966
		}, Vertex{
			x: -3.618034
			y: 0.0
			z: -1.381966
		}, Vertex{
			x: 1.381966
			y: 3.618034
			z: 0.0
		}, Vertex{
			x: 1.381966
			y: -3.618034
			z: 0.0
		}, Vertex{
			x: -1.381966
			y: 3.618034
			z: 0.0
		}, Vertex{
			x: -1.381966
			y: -3.618034
			z: 0.0
		}, Vertex{
			x: 2.170821
			y: 0.0
			z: 3.512461
		}, Vertex{
			x: 2.170821
			y: 0.0
			z: -3.512461
		}, Vertex{
			x: -2.170821
			y: 0.0
			z: 3.512461
		}, Vertex{
			x: -2.170821
			y: 0.0
			z: -3.512461
		}, Vertex{
			x: 3.512461
			y: 2.170821
			z: 0.0
		}, Vertex{
			x: 3.512461
			y: -2.170821
			z: 0.0
		}, Vertex{
			x: -3.512461
			y: 2.170821
			z: 0.0
		}, Vertex{
			x: -3.512461
			y: -2.170821
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 3.512461
			z: 2.170821
		}, Vertex{
			x: 0.0
			y: 3.512461
			z: -2.170821
		}, Vertex{
			x: 0.0
			y: -3.512461
			z: 2.170821
		}, Vertex{
			x: 0.0
			y: -3.512461
			z: -2.170821
		}, Vertex{
			x: 1.175186
			y: 1.901492
			z: 3.076678
		}, Vertex{
			x: 1.175186
			y: 1.901492
			z: -3.076678
		}, Vertex{
			x: 1.175186
			y: -1.901492
			z: 3.076678
		}, Vertex{
			x: 1.175186
			y: -1.901492
			z: -3.076678
		}, Vertex{
			x: -1.175186
			y: 1.901492
			z: 3.076678
		}, Vertex{
			x: -1.175186
			y: 1.901492
			z: -3.076678
		}, Vertex{
			x: -1.175186
			y: -1.901492
			z: 3.076678
		}, Vertex{
			x: -1.175186
			y: -1.901492
			z: -3.076678
		}, Vertex{
			x: 3.076678
			y: 1.175186
			z: 1.901492
		}, Vertex{
			x: 3.076678
			y: 1.175186
			z: -1.901492
		}, Vertex{
			x: 3.076678
			y: -1.175186
			z: 1.901492
		}, Vertex{
			x: 3.076678
			y: -1.175186
			z: -1.901492
		}, Vertex{
			x: -3.076678
			y: 1.175186
			z: 1.901492
		}, Vertex{
			x: -3.076678
			y: 1.175186
			z: -1.901492
		}, Vertex{
			x: -3.076678
			y: -1.175186
			z: 1.901492
		}, Vertex{
			x: -3.076678
			y: -1.175186
			z: -1.901492
		}, Vertex{
			x: 1.901492
			y: 3.076678
			z: 1.175186
		}, Vertex{
			x: 1.901492
			y: 3.076678
			z: -1.175186
		}, Vertex{
			x: 1.901492
			y: -3.076678
			z: 1.175186
		}, Vertex{
			x: 1.901492
			y: -3.076678
			z: -1.175186
		}, Vertex{
			x: -1.901492
			y: 3.076678
			z: 1.175186
		}, Vertex{
			x: -1.901492
			y: 3.076678
			z: -1.175186
		}, Vertex{
			x: -1.901492
			y: -3.076678
			z: 1.175186
		}, Vertex{
			x: -1.901492
			y: -3.076678
			z: -1.175186
		}, Vertex{
			x: 2.236068
			y: 2.236068
			z: 2.236068
		}, Vertex{
			x: 2.236068
			y: 2.236068
			z: -2.236068
		}, Vertex{
			x: 2.236068
			y: -2.236068
			z: 2.236068
		}, Vertex{
			x: 2.236068
			y: -2.236068
			z: -2.236068
		}, Vertex{
			x: -2.236068
			y: 2.236068
			z: 2.236068
		}, Vertex{
			x: -2.236068
			y: 2.236068
			z: -2.236068
		}, Vertex{
			x: -2.236068
			y: -2.236068
			z: 2.236068
		}, Vertex{
			x: -2.236068
			y: -2.236068
			z: -2.236068
		}]
		faces:     [[18, 0, 8], [18, 8, 32], [18, 32, 56], [18, 56, 40],
			[18, 40, 10], [18, 10, 38], [18, 38, 54], [18, 54, 30],
			[18, 30, 6], [18, 6, 0], [19, 1, 7], [19, 7, 31],
			[19, 31, 55], [19, 55, 39], [19, 39, 11], [19, 11, 41],
			[19, 41, 57], [19, 57, 33], [19, 33, 9], [19, 9, 1],
			[20, 0, 6], [20, 6, 34], [20, 34, 58], [20, 58, 42],
			[20, 42, 12], [20, 12, 44], [20, 44, 60], [20, 60, 36],
			[20, 36, 8], [20, 8, 0], [21, 1, 9], [21, 9, 37],
			[21, 37, 61], [21, 61, 45], [21, 45, 13], [21, 13, 43],
			[21, 43, 59], [21, 59, 35], [21, 35, 7], [21, 7, 1],
			[22, 2, 11], [22, 11, 39], [22, 39, 55], [22, 55, 47],
			[22, 47, 14], [22, 14, 46], [22, 46, 54], [22, 54, 38],
			[22, 38, 10], [22, 10, 2], [23, 2, 10], [23, 10, 40],
			[23, 40, 56], [23, 56, 48], [23, 48, 15], [23, 15, 49],
			[23, 49, 57], [23, 57, 41], [23, 41, 11], [23, 11, 2],
			[24, 3, 12], [24, 12, 42], [24, 42, 58], [24, 58, 50],
			[24, 50, 16], [24, 16, 51], [24, 51, 59], [24, 59, 43],
			[24, 43, 13], [24, 13, 3], [25, 3, 13], [25, 13, 45],
			[25, 45, 61], [25, 61, 53], [25, 53, 17], [25, 17, 52],
			[25, 52, 60], [25, 60, 44], [25, 44, 12], [25, 12, 3],
			[26, 4, 16], [26, 16, 50], [26, 50, 58], [26, 58, 34],
			[26, 34, 6], [26, 6, 30], [26, 30, 54], [26, 54, 46],
			[26, 46, 14], [26, 14, 4], [27, 4, 14], [27, 14, 47],
			[27, 47, 55], [27, 55, 31], [27, 31, 7], [27, 7, 35],
			[27, 35, 59], [27, 59, 51], [27, 51, 16], [27, 16, 4],
			[28, 5, 15], [28, 15, 48], [28, 48, 56], [28, 56, 32],
			[28, 32, 8], [28, 8, 36], [28, 36, 60], [28, 60, 52],
			[28, 52, 17], [28, 17, 5], [29, 5, 17], [29, 17, 53],
			[29, 53, 61], [29, 61, 37], [29, 37, 9], [29, 9, 33],
			[29, 33, 57], [29, 57, 49], [29, 49, 15], [29, 15, 5]]
	},
	Polyhedron{
		name:      'IcositruncatedDodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.1909830
			z: 1.927051
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: -1.927051
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: 1.927051
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: -1.927051
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: 1.927051
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: -1.927051
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: 1.927051
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: -1.927051
		}, Vertex{
			x: 1.927051
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: 1.927051
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: 1.927051
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: 1.927051
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: -1.927051
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -1.927051
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: -1.927051
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: -1.927051
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: 0.1909830
			y: 1.927051
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: 1.927051
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: -1.927051
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: -1.927051
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: 1.927051
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: 1.927051
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: -1.927051
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: -1.927051
			z: -0.5
		}, Vertex{
			x: 0.690983
			y: 0.5
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: 0.5
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: -0.5
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: -0.5
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: 0.5
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: 0.5
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: -0.5
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: -0.5
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: 0.5
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: -0.5
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: 0.5
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: -0.5
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: 0.5
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: -0.5
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: 0.5
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: 0.5
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: 0.5
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: 0.5
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: -0.5
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: -0.5
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: -0.5
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: -0.5
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: 1.0
			y: 0.618034
			z: 1.618034
		}, Vertex{
			x: 1.0
			y: 0.618034
			z: -1.618034
		}, Vertex{
			x: 1.0
			y: -0.618034
			z: 1.618034
		}, Vertex{
			x: 1.0
			y: -0.618034
			z: -1.618034
		}, Vertex{
			x: -1.0
			y: 0.618034
			z: 1.618034
		}, Vertex{
			x: -1.0
			y: 0.618034
			z: -1.618034
		}, Vertex{
			x: -1.0
			y: -0.618034
			z: 1.618034
		}, Vertex{
			x: -1.0
			y: -0.618034
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 1.0
			z: 0.618034
		}, Vertex{
			x: 1.618034
			y: 1.0
			z: -0.618034
		}, Vertex{
			x: 1.618034
			y: -1.0
			z: 0.618034
		}, Vertex{
			x: 1.618034
			y: -1.0
			z: -0.618034
		}, Vertex{
			x: -1.618034
			y: 1.0
			z: 0.618034
		}, Vertex{
			x: -1.618034
			y: 1.0
			z: -0.618034
		}, Vertex{
			x: -1.618034
			y: -1.0
			z: 0.618034
		}, Vertex{
			x: -1.618034
			y: -1.0
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 1.618034
			z: 1.0
		}, Vertex{
			x: 0.618034
			y: 1.618034
			z: -1.0
		}, Vertex{
			x: 0.618034
			y: -1.618034
			z: 1.0
		}, Vertex{
			x: 0.618034
			y: -1.618034
			z: -1.0
		}, Vertex{
			x: -0.618034
			y: 1.618034
			z: 1.0
		}, Vertex{
			x: -0.618034
			y: 1.618034
			z: -1.0
		}, Vertex{
			x: -0.618034
			y: -1.618034
			z: 1.0
		}, Vertex{
			x: -0.618034
			y: -1.618034
			z: -1.0
		}, Vertex{
			x: 0.1909830
			y: 1.309017
			z: 1.5
		}, Vertex{
			x: 0.1909830
			y: 1.309017
			z: -1.5
		}, Vertex{
			x: 0.1909830
			y: -1.309017
			z: 1.5
		}, Vertex{
			x: 0.1909830
			y: -1.309017
			z: -1.5
		}, Vertex{
			x: -0.1909830
			y: 1.309017
			z: 1.5
		}, Vertex{
			x: -0.1909830
			y: 1.309017
			z: -1.5
		}, Vertex{
			x: -0.1909830
			y: -1.309017
			z: 1.5
		}, Vertex{
			x: -0.1909830
			y: -1.309017
			z: -1.5
		}, Vertex{
			x: 1.5
			y: 0.1909830
			z: 1.309017
		}, Vertex{
			x: 1.5
			y: 0.1909830
			z: -1.309017
		}, Vertex{
			x: 1.5
			y: -0.1909830
			z: 1.309017
		}, Vertex{
			x: 1.5
			y: -0.1909830
			z: -1.309017
		}, Vertex{
			x: -1.5
			y: 0.1909830
			z: 1.309017
		}, Vertex{
			x: -1.5
			y: 0.1909830
			z: -1.309017
		}, Vertex{
			x: -1.5
			y: -0.1909830
			z: 1.309017
		}, Vertex{
			x: -1.5
			y: -0.1909830
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.5
			z: 0.1909830
		}, Vertex{
			x: 1.309017
			y: 1.5
			z: -0.1909830
		}, Vertex{
			x: 1.309017
			y: -1.5
			z: 0.1909830
		}, Vertex{
			x: 1.309017
			y: -1.5
			z: -0.1909830
		}, Vertex{
			x: -1.309017
			y: 1.5
			z: 0.1909830
		}, Vertex{
			x: -1.309017
			y: 1.5
			z: -0.1909830
		}, Vertex{
			x: -1.309017
			y: -1.5
			z: 0.1909830
		}, Vertex{
			x: -1.309017
			y: -1.5
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: 1.427051
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: 1.427051
			z: -1.309017
		}, Vertex{
			x: 0.5
			y: -1.427051
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: -1.427051
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: 1.427051
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: 1.427051
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: -1.427051
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: -1.427051
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: 1.427051
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: -1.427051
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: 1.427051
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: -1.427051
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: 1.427051
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: -1.427051
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: 1.427051
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: -1.427051
		}, Vertex{
			x: 1.427051
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: 1.427051
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: 1.427051
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: 1.427051
			y: -1.309017
			z: -0.5
		}, Vertex{
			x: -1.427051
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: -1.427051
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: -1.427051
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: -1.427051
			y: -1.309017
			z: -0.5
		}]
		faces:     [[0, 50, 80, 24, 26, 82, 48, 2, 106, 104],
			[1, 105, 107, 3, 49, 83, 27, 25, 81, 51], [4, 108, 110, 6, 52, 86, 30, 28, 84, 54],
			[5, 55, 85, 29, 31, 87, 53, 7, 111, 109], [8, 57, 88, 32, 33, 89, 56, 9, 113, 112],
			[10, 114, 115, 11, 58, 91, 35, 34, 90, 59], [12, 116, 117, 13, 60, 93, 37, 36, 92, 61],
			[14, 63, 94, 38, 39, 95, 62, 15, 119, 118], [16, 68, 72, 40, 44, 76, 64, 20, 100, 96],
			[17, 97, 101, 21, 65, 77, 45, 41, 73, 69], [18, 98, 102, 22, 66, 78, 46, 42, 74, 70],
			[19, 71, 75, 43, 47, 79, 67, 23, 103, 99], [0, 104, 56, 89, 41, 45, 93, 60, 108, 4],
			[1, 5, 109, 61, 92, 44, 40, 88, 57, 105], [2, 6, 110, 62, 95, 47, 43, 91, 58, 106],
			[3, 107, 59, 90, 42, 46, 94, 63, 111, 7], [8, 112, 64, 76, 28, 30, 78, 66, 114, 10],
			[9, 11, 115, 67, 79, 31, 29, 77, 65, 113], [12, 14, 118, 70, 74, 26, 24, 72, 68, 116],
			[13, 117, 69, 73, 25, 27, 75, 71, 119, 15], [16, 96, 48, 82, 34, 35, 83, 49, 97, 17],
			[18, 19, 99, 51, 81, 33, 32, 80, 50, 98], [20, 21, 101, 53, 87, 39, 38, 86, 52, 100],
			[22, 102, 54, 84, 36, 37, 85, 55, 103, 23], [0, 4, 54, 102, 98, 50],
			[1, 51, 99, 103, 55, 5], [2, 48, 96, 100, 52, 6],
			[3, 7, 53, 101, 97, 49], [8, 10, 59, 107, 105, 57],
			[9, 56, 104, 106, 58, 11], [12, 61, 109, 111, 63, 14],
			[13, 15, 62, 110, 108, 60], [16, 17, 69, 117, 116, 68],
			[18, 70, 118, 119, 71, 19], [20, 64, 112, 113, 65, 21],
			[22, 23, 67, 115, 114, 66], [24, 80, 32, 88, 40, 72],
			[25, 73, 41, 89, 33, 81], [26, 74, 42, 90, 34, 82],
			[27, 83, 35, 91, 43, 75], [28, 76, 44, 92, 36, 84],
			[29, 85, 37, 93, 45, 77], [30, 86, 38, 94, 46, 78],
			[31, 79, 47, 95, 39, 87]]
	},
	Polyhedron{
		name:      'SmallDitrigonalDodecicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.309017
			z: 1.618034
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: -1.618034
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: 1.618034
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: -1.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: 1.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: -1.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: 1.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: 1.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: 1.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 1.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: -1.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: -1.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: -1.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: -1.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: 1.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: 1.618034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: -1.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: -1.618034
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: 1.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: 1.618034
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: -1.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: -1.618034
			z: -0.5
		}, Vertex{
			x: 0.0
			y: 1.118034
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 1.118034
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -1.118034
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -1.118034
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 1.118034
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -1.118034
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 1.118034
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 1.118034
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 1.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 1.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 1.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: -1.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: -1.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: -1.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: -1.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 1.0
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: -1.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: -1.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 1.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 1.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: -1.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: -1.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 1.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: -1.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 1.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: -1.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 1.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: -1.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 1.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: -1.0
		}]
		faces:     [[0, 4, 30, 14, 51, 59, 55, 47, 10, 28], [0, 38, 46, 47, 39, 1, 25, 21, 20, 24],
			[2, 26, 22, 23, 27, 3, 37, 45, 44, 36], [2, 28, 8, 45, 53, 57, 49, 12, 30, 6],
			[5, 1, 29, 11, 46, 54, 58, 50, 15, 31], [5, 43, 51, 50, 42, 4, 24, 16, 17, 25],
			[7, 27, 19, 18, 26, 6, 40, 48, 49, 41], [7, 31, 13, 48, 56, 52, 44, 9, 29, 3],
			[33, 11, 9, 32, 16, 56, 40, 42, 58, 18], [33, 19, 59, 43, 41, 57, 17, 32, 8, 10],
			[34, 13, 15, 35, 22, 54, 38, 36, 52, 20], [34, 21, 53, 37, 39, 55, 23, 35, 14, 12],
			[24, 20, 52, 56, 16], [25, 17, 57, 53, 21], [26, 18, 58, 54, 22],
			[27, 23, 55, 59, 19], [28, 2, 36, 38, 0], [29, 1, 39, 37, 3],
			[30, 4, 42, 40, 6], [31, 7, 41, 43, 5], [32, 9, 44, 45, 8],
			[33, 10, 47, 46, 11], [34, 12, 49, 48, 13], [35, 15, 50, 51, 14],
			[24, 4, 0], [25, 1, 5], [26, 2, 6], [27, 7, 3], [28, 10, 8],
			[29, 9, 11], [30, 12, 14], [31, 15, 13], [32, 17, 16],
			[33, 18, 19], [34, 20, 21], [35, 23, 22], [36, 44, 52],
			[37, 53, 45], [38, 54, 46], [39, 47, 55], [40, 56, 48],
			[41, 49, 57], [42, 50, 58], [43, 59, 51]]
	},
	Polyhedron{
		name:      'Rhombicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: 2.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 2.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: -0.5
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: 1.618034
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: -1.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: 1.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: -1.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: 1.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: -1.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: 1.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: 1.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: 1.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: 1.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: -1.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: -1.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: -1.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: -1.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: 1.618034
			z: -1.309017
		}, Vertex{
			x: 0.809017
			y: -1.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: -1.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: 1.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: 1.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: -1.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: -1.618034
			z: -1.309017
		}]
		faces:     [[24, 52, 16, 20, 56], [25, 57, 21, 17, 53],
			[26, 58, 22, 18, 54], [27, 55, 19, 23, 59], [28, 36, 0, 2, 38],
			[29, 39, 3, 1, 37], [30, 42, 6, 4, 40], [31, 41, 5, 7, 43],
			[32, 44, 8, 9, 45], [33, 47, 11, 10, 46], [34, 49, 13, 12, 48],
			[35, 50, 14, 15, 51], [0, 36, 52, 24], [1, 25, 53, 37],
			[2, 26, 54, 38], [3, 39, 55, 27], [4, 24, 56, 40],
			[5, 41, 57, 25], [6, 42, 58, 26], [7, 27, 59, 43],
			[8, 44, 36, 28], [9, 29, 37, 45], [10, 28, 38, 46],
			[11, 47, 39, 29], [12, 30, 40, 48], [13, 49, 41, 31],
			[14, 50, 42, 30], [15, 31, 43, 51], [16, 52, 44, 32],
			[17, 32, 45, 53], [18, 33, 46, 54], [19, 55, 47, 33],
			[20, 34, 48, 56], [21, 57, 49, 34], [22, 58, 50, 35],
			[23, 35, 51, 59], [0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9],
			[12, 13, 15, 14], [16, 17, 21, 20], [18, 22, 23, 19],
			[24, 4, 0], [25, 1, 5], [26, 2, 6], [27, 7, 3], [28, 10, 8],
			[29, 9, 11], [30, 12, 14], [31, 15, 13], [32, 17, 16],
			[33, 18, 19], [34, 20, 21], [35, 23, 22], [36, 44, 52],
			[37, 53, 45], [38, 54, 46], [39, 47, 55], [40, 56, 48],
			[41, 49, 57], [42, 50, 58], [43, 59, 51]]
	},
	Polyhedron{
		name:      'GreatTriambicIcosahedron'
		vertexes_: [Vertex{
			x: 0.7236068
			y: 0.0
			z: 0.2763932
		}, Vertex{
			x: 0.7236068
			y: 0.0
			z: -0.2763932
		}, Vertex{
			x: -0.7236068
			y: 0.0
			z: 0.2763932
		}, Vertex{
			x: -0.7236068
			y: 0.0
			z: -0.2763932
		}, Vertex{
			x: 0.0
			y: 0.2763932
			z: 0.7236068
		}, Vertex{
			x: 0.0
			y: 0.2763932
			z: -0.7236068
		}, Vertex{
			x: 0.0
			y: -0.2763932
			z: 0.7236068
		}, Vertex{
			x: 0.0
			y: -0.2763932
			z: -0.7236068
		}, Vertex{
			x: 0.2763932
			y: 0.7236068
			z: 0.0
		}, Vertex{
			x: -0.2763932
			y: 0.7236068
			z: 0.0
		}, Vertex{
			x: 0.2763932
			y: -0.7236068
			z: 0.0
		}, Vertex{
			x: -0.2763932
			y: -0.7236068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: 1.618034
		}, Vertex{
			x: 2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: -0.4472136
			y: -0.4472136
			z: -0.4472136
		}, Vertex{
			x: -0.4472136
			y: -0.4472136
			z: 0.4472136
		}, Vertex{
			x: 0.4472136
			y: -0.4472136
			z: -0.4472136
		}, Vertex{
			x: 0.4472136
			y: -0.4472136
			z: 0.4472136
		}, Vertex{
			x: -0.4472136
			y: 0.4472136
			z: -0.4472136
		}, Vertex{
			x: -0.4472136
			y: 0.4472136
			z: 0.4472136
		}, Vertex{
			x: 0.4472136
			y: 0.4472136
			z: -0.4472136
		}, Vertex{
			x: 0.4472136
			y: 0.4472136
			z: 0.4472136
		}]
		faces:     [[12, 0, 14, 30, 22, 26], [12, 26, 17, 5, 16, 24],
			[12, 24, 20, 28, 14, 2], [12, 2, 22, 9, 17, 4], [12, 4, 16, 8, 20, 0],
			[15, 1, 13, 27, 23, 31], [15, 31, 19, 6, 18, 29],
			[15, 29, 21, 25, 13, 3], [15, 3, 23, 11, 19, 7], [15, 7, 18, 10, 21, 1],
			[13, 1, 21, 8, 16, 5], [13, 5, 17, 9, 23, 3], [13, 25, 16, 4, 17, 27],
			[14, 0, 20, 10, 18, 6], [14, 6, 19, 11, 22, 2], [14, 28, 18, 7, 19, 30],
			[20, 8, 21, 29, 18, 28], [20, 24, 16, 25, 21, 10],
			[22, 11, 23, 27, 17, 26], [22, 30, 19, 31, 23, 9]]
	},
	Polyhedron{
		name:      'GreatRhombicTriacontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: -0.3454915
			z: 0.2135255
		}, Vertex{
			x: 0.0
			y: -0.3454915
			z: -0.2135255
		}, Vertex{
			x: 0.0
			y: 0.3454915
			z: 0.2135255
		}, Vertex{
			x: 0.0
			y: 0.3454915
			z: -0.2135255
		}, Vertex{
			x: -0.3454915
			y: 0.2135255
			z: 0.0
		}, Vertex{
			x: 0.3454915
			y: 0.2135255
			z: 0.0
		}, Vertex{
			x: -0.3454915
			y: -0.2135255
			z: 0.0
		}, Vertex{
			x: 0.3454915
			y: -0.2135255
			z: 0.0
		}, Vertex{
			x: 0.2135255
			y: 0.0
			z: -0.3454915
		}, Vertex{
			x: 0.2135255
			y: 0.0
			z: 0.3454915
		}, Vertex{
			x: -0.2135255
			y: 0.0
			z: -0.3454915
		}, Vertex{
			x: -0.2135255
			y: 0.0
			z: 0.3454915
		}, Vertex{
			x: 0.559017
			y: 0.0
			z: 0.2135255
		}, Vertex{
			x: 0.559017
			y: 0.0
			z: -0.2135255
		}, Vertex{
			x: -0.559017
			y: 0.0
			z: 0.2135255
		}, Vertex{
			x: -0.559017
			y: 0.0
			z: -0.2135255
		}, Vertex{
			x: 0.0
			y: 0.2135255
			z: 0.559017
		}, Vertex{
			x: 0.0
			y: 0.2135255
			z: -0.559017
		}, Vertex{
			x: 0.0
			y: -0.2135255
			z: 0.559017
		}, Vertex{
			x: 0.0
			y: -0.2135255
			z: -0.559017
		}, Vertex{
			x: 0.2135255
			y: 0.559017
			z: 0.0
		}, Vertex{
			x: -0.2135255
			y: 0.559017
			z: 0.0
		}, Vertex{
			x: 0.2135255
			y: -0.559017
			z: 0.0
		}, Vertex{
			x: -0.2135255
			y: -0.559017
			z: 0.0
		}, Vertex{
			x: -0.3454915
			y: -0.3454915
			z: -0.3454915
		}, Vertex{
			x: -0.3454915
			y: -0.3454915
			z: 0.3454915
		}, Vertex{
			x: 0.3454915
			y: -0.3454915
			z: -0.3454915
		}, Vertex{
			x: 0.3454915
			y: -0.3454915
			z: 0.3454915
		}, Vertex{
			x: -0.3454915
			y: 0.3454915
			z: -0.3454915
		}, Vertex{
			x: -0.3454915
			y: 0.3454915
			z: 0.3454915
		}, Vertex{
			x: 0.3454915
			y: 0.3454915
			z: -0.3454915
		}, Vertex{
			x: 0.3454915
			y: 0.3454915
			z: 0.3454915
		}]
		faces:     [[0, 12, 2, 14], [0, 14, 10, 26], [0, 26, 5, 16],
			[1, 13, 9, 25], [1, 25, 4, 17], [1, 17, 5, 27], [2, 28, 6, 18],
			[2, 18, 7, 30], [2, 30, 10, 14], [3, 19, 6, 29], [3, 29, 9, 13],
			[3, 13, 1, 15], [4, 20, 8, 24], [4, 24, 0, 16], [4, 16, 5, 17],
			[7, 18, 6, 19], [7, 19, 3, 31], [7, 31, 11, 23], [8, 22, 6, 28],
			[8, 28, 2, 12], [8, 12, 0, 24], [9, 29, 6, 22], [9, 22, 8, 20],
			[9, 20, 4, 25], [10, 30, 7, 23], [10, 23, 11, 21],
			[10, 21, 5, 26], [11, 31, 3, 15], [11, 15, 1, 27],
			[11, 27, 5, 21]]
	},
	Polyhedron{
		name:      'GreatHexagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.1717804
			y: 0.05943847
			z: 0.5847722
		}, Vertex{
			x: 0.1717804
			y: -0.05943847
			z: -0.5847722
		}, Vertex{
			x: -0.1717804
			y: -0.05943847
			z: 0.5847722
		}, Vertex{
			x: -0.1717804
			y: 0.05943847
			z: -0.5847722
		}, Vertex{
			x: 0.5847722
			y: 0.1717804
			z: 0.05943847
		}, Vertex{
			x: 0.5847722
			y: -0.1717804
			z: -0.05943847
		}, Vertex{
			x: -0.5847722
			y: -0.1717804
			z: 0.05943847
		}, Vertex{
			x: -0.5847722
			y: 0.1717804
			z: -0.05943847
		}, Vertex{
			x: 0.05943847
			y: 0.5847722
			z: 0.1717804
		}, Vertex{
			x: 0.05943847
			y: -0.5847722
			z: -0.1717804
		}, Vertex{
			x: -0.05943847
			y: -0.5847722
			z: 0.1717804
		}, Vertex{
			x: -0.05943847
			y: 0.5847722
			z: -0.1717804
		}, Vertex{
			x: 0.0
			y: 0.218508
			z: 0.5720614
		}, Vertex{
			x: 0.0
			y: 0.218508
			z: -0.5720614
		}, Vertex{
			x: 0.0
			y: -0.218508
			z: 0.5720614
		}, Vertex{
			x: 0.0
			y: -0.218508
			z: -0.5720614
		}, Vertex{
			x: 0.5720614
			y: 0.0
			z: 0.218508
		}, Vertex{
			x: 0.5720614
			y: 0.0
			z: -0.218508
		}, Vertex{
			x: -0.5720614
			y: 0.0
			z: 0.218508
		}, Vertex{
			x: -0.5720614
			y: 0.0
			z: -0.218508
		}, Vertex{
			x: 0.218508
			y: 0.5720614
			z: 0.0
		}, Vertex{
			x: 0.218508
			y: -0.5720614
			z: 0.0
		}, Vertex{
			x: -0.218508
			y: 0.5720614
			z: 0.0
		}, Vertex{
			x: -0.218508
			y: -0.5720614
			z: 0.0
		}, Vertex{
			x: 0.218508
			y: -0.1350454
			z: 0.5558929
		}, Vertex{
			x: 0.218508
			y: 0.1350454
			z: -0.5558929
		}, Vertex{
			x: -0.218508
			y: 0.1350454
			z: 0.5558929
		}, Vertex{
			x: -0.218508
			y: -0.1350454
			z: -0.5558929
		}, Vertex{
			x: 0.5558929
			y: -0.218508
			z: 0.1350454
		}, Vertex{
			x: 0.5558929
			y: 0.218508
			z: -0.1350454
		}, Vertex{
			x: -0.5558929
			y: 0.218508
			z: 0.1350454
		}, Vertex{
			x: -0.5558929
			y: -0.218508
			z: -0.1350454
		}, Vertex{
			x: 0.1350454
			y: -0.5558929
			z: 0.218508
		}, Vertex{
			x: 0.1350454
			y: 0.5558929
			z: -0.218508
		}, Vertex{
			x: -0.1350454
			y: 0.5558929
			z: 0.218508
		}, Vertex{
			x: -0.1350454
			y: -0.5558929
			z: -0.218508
		}, Vertex{
			x: 0.3146815
			y: 0.1717804
			z: 0.4964545
		}, Vertex{
			x: 0.3146815
			y: -0.1717804
			z: -0.4964545
		}, Vertex{
			x: -0.3146815
			y: -0.1717804
			z: 0.4964545
		}, Vertex{
			x: -0.3146815
			y: 0.1717804
			z: -0.4964545
		}, Vertex{
			x: 0.4964545
			y: 0.3146815
			z: 0.1717804
		}, Vertex{
			x: 0.4964545
			y: -0.3146815
			z: -0.1717804
		}, Vertex{
			x: -0.4964545
			y: -0.3146815
			z: 0.1717804
		}, Vertex{
			x: -0.4964545
			y: 0.3146815
			z: -0.1717804
		}, Vertex{
			x: 0.1717804
			y: 0.4964545
			z: 0.3146815
		}, Vertex{
			x: 0.1717804
			y: -0.4964545
			z: -0.3146815
		}, Vertex{
			x: -0.1717804
			y: -0.4964545
			z: 0.3146815
		}, Vertex{
			x: -0.1717804
			y: 0.4964545
			z: -0.3146815
		}, Vertex{
			x: 0.2779465
			y: 0.0
			z: 0.4497269
		}, Vertex{
			x: 0.2779465
			y: 0.0
			z: 0.4497269
		}, Vertex{
			x: 0.2779465
			y: 0.0
			z: -0.4497269
		}, Vertex{
			x: 0.2779465
			y: 0.0
			z: -0.4497269
		}, Vertex{
			x: -0.2779465
			y: 0.0
			z: 0.4497269
		}, Vertex{
			x: -0.2779465
			y: 0.0
			z: 0.4497269
		}, Vertex{
			x: -0.2779465
			y: 0.0
			z: -0.4497269
		}, Vertex{
			x: -0.2779465
			y: 0.0
			z: -0.4497269
		}, Vertex{
			x: 0.4497269
			y: 0.2779465
			z: 0.0
		}, Vertex{
			x: 0.4497269
			y: 0.2779465
			z: 0.0
		}, Vertex{
			x: 0.4497269
			y: -0.2779465
			z: 0.0
		}, Vertex{
			x: 0.4497269
			y: -0.2779465
			z: 0.0
		}, Vertex{
			x: -0.4497269
			y: 0.2779465
			z: 0.0
		}, Vertex{
			x: -0.4497269
			y: 0.2779465
			z: 0.0
		}, Vertex{
			x: -0.4497269
			y: -0.2779465
			z: 0.0
		}, Vertex{
			x: -0.4497269
			y: -0.2779465
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.4497269
			z: 0.2779465
		}, Vertex{
			x: 0.0
			y: 0.4497269
			z: 0.2779465
		}, Vertex{
			x: 0.0
			y: 0.4497269
			z: -0.2779465
		}, Vertex{
			x: 0.0
			y: 0.4497269
			z: -0.2779465
		}, Vertex{
			x: 0.0
			y: -0.4497269
			z: 0.2779465
		}, Vertex{
			x: 0.0
			y: -0.4497269
			z: 0.2779465
		}, Vertex{
			x: 0.0
			y: -0.4497269
			z: -0.2779465
		}, Vertex{
			x: 0.0
			y: -0.4497269
			z: -0.2779465
		}, Vertex{
			x: 0.3902884
			y: -0.1429011
			z: 0.4497269
		}, Vertex{
			x: 0.3902884
			y: 0.1429011
			z: -0.4497269
		}, Vertex{
			x: -0.3902884
			y: 0.1429011
			z: 0.4497269
		}, Vertex{
			x: -0.3902884
			y: -0.1429011
			z: -0.4497269
		}, Vertex{
			x: 0.4497269
			y: -0.3902884
			z: 0.1429011
		}, Vertex{
			x: 0.4497269
			y: 0.3902884
			z: -0.1429011
		}, Vertex{
			x: -0.4497269
			y: 0.3902884
			z: 0.1429011
		}, Vertex{
			x: -0.4497269
			y: -0.3902884
			z: -0.1429011
		}, Vertex{
			x: 0.1429011
			y: -0.4497269
			z: 0.3902884
		}, Vertex{
			x: 0.1429011
			y: 0.4497269
			z: -0.3902884
		}, Vertex{
			x: -0.1429011
			y: 0.4497269
			z: 0.3902884
		}, Vertex{
			x: -0.1429011
			y: -0.4497269
			z: -0.3902884
		}, Vertex{
			x: 0.04672764
			y: 0.4129919
			z: 0.4497269
		}, Vertex{
			x: 0.04672764
			y: -0.4129919
			z: -0.4497269
		}, Vertex{
			x: -0.04672764
			y: -0.4129919
			z: 0.4497269
		}, Vertex{
			x: -0.04672764
			y: 0.4129919
			z: -0.4497269
		}, Vertex{
			x: 0.4497269
			y: 0.04672764
			z: 0.4129919
		}, Vertex{
			x: 0.4497269
			y: -0.04672764
			z: -0.4129919
		}, Vertex{
			x: -0.4497269
			y: -0.04672764
			z: 0.4129919
		}, Vertex{
			x: -0.4497269
			y: 0.04672764
			z: -0.4129919
		}, Vertex{
			x: 0.4129919
			y: 0.4497269
			z: 0.04672764
		}, Vertex{
			x: 0.4129919
			y: -0.4497269
			z: -0.04672764
		}, Vertex{
			x: -0.4129919
			y: -0.4497269
			z: 0.04672764
		}, Vertex{
			x: -0.4129919
			y: 0.4497269
			z: -0.04672764
		}, Vertex{
			x: 0.3535534
			y: 0.3535534
			z: 0.3535534
		}, Vertex{
			x: 0.3535534
			y: 0.3535534
			z: -0.3535534
		}, Vertex{
			x: 0.3535534
			y: -0.3535534
			z: 0.3535534
		}, Vertex{
			x: 0.3535534
			y: -0.3535534
			z: -0.3535534
		}, Vertex{
			x: -0.3535534
			y: 0.3535534
			z: 0.3535534
		}, Vertex{
			x: -0.3535534
			y: 0.3535534
			z: -0.3535534
		}, Vertex{
			x: -0.3535534
			y: -0.3535534
			z: 0.3535534
		}, Vertex{
			x: -0.3535534
			y: -0.3535534
			z: -0.3535534
		}]
		faces:     [[12, 30, 62, 10, 68, 80], [12, 80, 59, 29, 57, 92],
			[12, 92, 67, 43, 60, 30], [13, 29, 59, 9, 71, 83],
			[13, 83, 62, 30, 60, 95], [13, 95, 64, 40, 57, 29],
			[14, 28, 56, 8, 65, 82], [14, 82, 61, 31, 63, 94],
			[14, 94, 70, 41, 58, 28], [15, 31, 61, 11, 66, 81],
			[15, 81, 56, 28, 58, 93], [15, 93, 69, 42, 63, 31],
			[16, 32, 70, 1, 51, 73], [16, 73, 67, 34, 65, 84],
			[16, 84, 52, 46, 68, 32], [17, 33, 64, 0, 48, 72],
			[17, 72, 69, 35, 71, 85], [17, 85, 55, 47, 66, 33],
			[18, 34, 67, 3, 54, 75], [18, 75, 70, 32, 68, 86],
			[18, 86, 49, 44, 65, 34], [19, 35, 69, 2, 53, 74],
			[19, 74, 64, 33, 66, 87], [19, 87, 50, 45, 71, 35],
			[20, 25, 55, 7, 60, 78], [20, 78, 52, 24, 48, 88],
			[20, 88, 59, 37, 51, 25], [21, 24, 52, 6, 63, 79],
			[21, 79, 55, 25, 51, 89], [21, 89, 56, 36, 48, 24],
			[22, 26, 49, 4, 57, 77], [22, 77, 50, 27, 54, 91],
			[22, 91, 62, 38, 53, 26], [23, 27, 50, 5, 58, 76],
			[23, 76, 49, 26, 53, 90], [23, 90, 61, 39, 54, 27],
			[96, 2, 69, 93, 58, 5], [96, 5, 50, 87, 66, 11], [96, 11, 61, 90, 53, 2],
			[97, 39, 61, 82, 65, 44], [97, 44, 49, 76, 58, 41],
			[97, 41, 70, 75, 54, 39], [98, 38, 62, 83, 71, 45],
			[98, 45, 50, 77, 57, 40], [98, 40, 64, 74, 53, 38],
			[99, 3, 67, 92, 57, 4], [99, 4, 49, 86, 68, 10], [99, 10, 62, 91, 54, 3],
			[100, 36, 56, 81, 66, 47], [100, 47, 55, 79, 63, 42],
			[100, 42, 69, 72, 48, 36], [101, 1, 70, 94, 63, 6],
			[101, 6, 52, 84, 65, 8], [101, 8, 56, 89, 51, 1],
			[102, 0, 64, 95, 60, 7], [102, 7, 55, 85, 71, 9],
			[102, 9, 59, 88, 48, 0], [103, 37, 59, 80, 68, 46],
			[103, 46, 52, 78, 60, 43], [103, 43, 67, 73, 51, 37]]
	},
	Polyhedron{
		name:      'SnubCube(laevo}'
		vertexes_: [Vertex{
			x: 0.6212264
			y: 0.3377540
			z: 1.142614
		}, Vertex{
			x: 0.6212264
			y: -0.3377540
			z: -1.142614
		}, Vertex{
			x: -0.6212264
			y: -0.3377540
			z: 1.142614
		}, Vertex{
			x: -0.6212264
			y: 0.3377540
			z: -1.142614
		}, Vertex{
			x: 1.142614
			y: 0.6212264
			z: 0.3377540
		}, Vertex{
			x: 1.142614
			y: -0.6212264
			z: -0.3377540
		}, Vertex{
			x: -1.142614
			y: -0.6212264
			z: 0.3377540
		}, Vertex{
			x: -1.142614
			y: 0.6212264
			z: -0.3377540
		}, Vertex{
			x: 0.3377540
			y: 1.142614
			z: 0.6212264
		}, Vertex{
			x: 0.3377540
			y: -1.142614
			z: -0.6212264
		}, Vertex{
			x: -0.3377540
			y: -1.142614
			z: 0.6212264
		}, Vertex{
			x: -0.3377540
			y: 1.142614
			z: -0.6212264
		}, Vertex{
			x: 0.3377540
			y: -0.6212264
			z: 1.142614
		}, Vertex{
			x: 0.3377540
			y: 0.6212264
			z: -1.142614
		}, Vertex{
			x: -0.3377540
			y: 0.6212264
			z: 1.142614
		}, Vertex{
			x: -0.3377540
			y: -0.6212264
			z: -1.142614
		}, Vertex{
			x: 1.142614
			y: -0.3377540
			z: 0.6212264
		}, Vertex{
			x: 1.142614
			y: 0.3377540
			z: -0.6212264
		}, Vertex{
			x: -1.142614
			y: 0.3377540
			z: 0.6212264
		}, Vertex{
			x: -1.142614
			y: -0.3377540
			z: -0.6212264
		}, Vertex{
			x: 0.6212264
			y: -1.142614
			z: 0.3377540
		}, Vertex{
			x: 0.6212264
			y: 1.142614
			z: -0.3377540
		}, Vertex{
			x: -0.6212264
			y: 1.142614
			z: 0.3377540
		}, Vertex{
			x: -0.6212264
			y: -1.142614
			z: -0.3377540
		}]
		faces:     [[2, 12, 0, 14], [3, 13, 1, 15], [4, 16, 5, 17],
			[7, 19, 6, 18], [8, 21, 11, 22], [9, 20, 10, 23],
			[0, 8, 14], [1, 9, 15], [2, 10, 12], [3, 11, 13],
			[4, 0, 16], [5, 1, 17], [6, 2, 18], [7, 3, 19], [8, 4, 21],
			[9, 5, 20], [10, 6, 23], [11, 7, 22], [12, 16, 0],
			[13, 17, 1], [14, 18, 2], [15, 19, 3], [16, 20, 5],
			[17, 21, 4], [18, 22, 7], [19, 23, 6], [20, 12, 10],
			[21, 13, 11], [22, 14, 8], [23, 15, 9], [8, 0, 4],
			[9, 1, 5], [10, 2, 6], [11, 3, 7], [12, 20, 16], [13, 21, 17],
			[14, 22, 18], [15, 23, 19]]
	},
	Polyhedron{
		name:      'TriakisOctahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 2.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -2.414214
		}, Vertex{
			x: 2.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -2.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -2.414214
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[6, 0, 2], [6, 2, 4], [6, 4, 0], [7, 1, 4],
			[7, 4, 2], [7, 2, 1], [8, 0, 5], [8, 5, 2], [8, 2, 0],
			[9, 1, 2], [9, 2, 5], [9, 5, 1], [10, 0, 4], [10, 4, 3],
			[10, 3, 0], [11, 1, 3], [11, 3, 4], [11, 4, 1], [12, 0, 3],
			[12, 3, 5], [12, 5, 0], [13, 1, 5], [13, 5, 3], [13, 3, 1]]
	},
	Polyhedron{
		name:      'PentagonalIcositetrahedron(dextro}'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.361410
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.361410
		}, Vertex{
			x: 1.361410
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.361410
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.361410
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.361410
			z: 0.0
		}, Vertex{
			x: 0.7401838
			y: -0.2187966
			z: 1.023656
		}, Vertex{
			x: 0.7401838
			y: 0.2187966
			z: -1.023656
		}, Vertex{
			x: -0.7401838
			y: 0.2187966
			z: 1.023656
		}, Vertex{
			x: -0.7401838
			y: -0.2187966
			z: -1.023656
		}, Vertex{
			x: 1.023656
			y: -0.7401838
			z: 0.2187966
		}, Vertex{
			x: 1.023656
			y: 0.7401838
			z: -0.2187966
		}, Vertex{
			x: -1.023656
			y: 0.7401838
			z: 0.2187966
		}, Vertex{
			x: -1.023656
			y: -0.7401838
			z: -0.2187966
		}, Vertex{
			x: 0.2187966
			y: -1.023656
			z: 0.7401838
		}, Vertex{
			x: 0.2187966
			y: 1.023656
			z: -0.7401838
		}, Vertex{
			x: -0.2187966
			y: 1.023656
			z: 0.7401838
		}, Vertex{
			x: -0.2187966
			y: -1.023656
			z: -0.7401838
		}, Vertex{
			x: 0.2187966
			y: 0.7401838
			z: 1.023656
		}, Vertex{
			x: 0.2187966
			y: -0.7401838
			z: -1.023656
		}, Vertex{
			x: -0.2187966
			y: -0.7401838
			z: 1.023656
		}, Vertex{
			x: -0.2187966
			y: 0.7401838
			z: -1.023656
		}, Vertex{
			x: 1.023656
			y: 0.2187966
			z: 0.7401838
		}, Vertex{
			x: 1.023656
			y: -0.2187966
			z: -0.7401838
		}, Vertex{
			x: -1.023656
			y: -0.2187966
			z: 0.7401838
		}, Vertex{
			x: -1.023656
			y: 0.2187966
			z: -0.7401838
		}, Vertex{
			x: 0.7401838
			y: 1.023656
			z: 0.2187966
		}, Vertex{
			x: 0.7401838
			y: -1.023656
			z: -0.2187966
		}, Vertex{
			x: -0.7401838
			y: -1.023656
			z: 0.2187966
		}, Vertex{
			x: -0.7401838
			y: 1.023656
			z: -0.2187966
		}, Vertex{
			x: 0.7401838
			y: 0.7401838
			z: 0.7401838
		}, Vertex{
			x: 0.7401838
			y: 0.7401838
			z: -0.7401838
		}, Vertex{
			x: 0.7401838
			y: -0.7401838
			z: 0.7401838
		}, Vertex{
			x: 0.7401838
			y: -0.7401838
			z: -0.7401838
		}, Vertex{
			x: -0.7401838
			y: 0.7401838
			z: 0.7401838
		}, Vertex{
			x: -0.7401838
			y: 0.7401838
			z: -0.7401838
		}, Vertex{
			x: -0.7401838
			y: -0.7401838
			z: 0.7401838
		}, Vertex{
			x: -0.7401838
			y: -0.7401838
			z: -0.7401838
		}]
		faces:     [[0, 6, 22, 30, 18], [0, 18, 16, 34, 8], [0, 8, 24, 36, 20],
			[0, 20, 14, 32, 6], [1, 7, 23, 33, 19], [1, 19, 17, 37, 9],
			[1, 9, 25, 35, 21], [1, 21, 15, 31, 7], [2, 10, 27, 33, 23],
			[2, 23, 7, 31, 11], [2, 11, 26, 30, 22], [2, 22, 6, 32, 10],
			[3, 12, 29, 35, 25], [3, 25, 9, 37, 13], [3, 13, 28, 36, 24],
			[3, 24, 8, 34, 12], [4, 15, 21, 35, 29], [4, 29, 12, 34, 16],
			[4, 16, 18, 30, 26], [4, 26, 11, 31, 15], [5, 14, 20, 36, 28],
			[5, 28, 13, 37, 17], [5, 17, 19, 33, 27], [5, 27, 10, 32, 14]]
	},
	Polyhedron{
		name:      'GreatDitrigonalIcosidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: 0.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: 0.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: 0.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: 0.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: 0.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: 0.0
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.5
		}]
		faces:     [[0, 6, 19, 15, 4], [0, 8, 1, 19, 18], [0, 14, 15, 1, 10],
			[7, 1, 5, 14, 18], [7, 11, 14, 12, 10], [7, 16, 12, 5, 3],
			[9, 2, 16, 17, 3], [9, 5, 8, 16, 18], [9, 19, 17, 8, 4],
			[13, 12, 2, 11, 3], [13, 15, 11, 6, 10], [13, 17, 6, 2, 4],
			[0, 4, 8], [0, 10, 6], [0, 18, 14], [1, 7, 10], [1, 8, 5],
			[1, 15, 19], [2, 6, 11], [2, 9, 4], [2, 12, 16], [3, 5, 9],
			[3, 11, 7], [3, 17, 13], [4, 15, 13], [5, 12, 14],
			[6, 17, 19], [7, 18, 16], [8, 17, 16], [9, 18, 19],
			[10, 12, 13], [11, 15, 14]]
	},
	Polyhedron{
		name:      'GreatDodecicosacron'
		vertexes_: [Vertex{
			x: 0.0
			y: -0.927051
			z: 0.572949
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: -0.572949
		}, Vertex{
			x: 0.0
			y: 0.927051
			z: 0.572949
		}, Vertex{
			x: 0.0
			y: 0.927051
			z: -0.572949
		}, Vertex{
			x: -0.927051
			y: 0.572949
			z: 0.0
		}, Vertex{
			x: 0.927051
			y: 0.572949
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: -0.572949
			z: 0.0
		}, Vertex{
			x: 0.927051
			y: -0.572949
			z: 0.0
		}, Vertex{
			x: 0.572949
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: 0.572949
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: -0.572949
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: -0.572949
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: 1.118034
		}]
		faces:     [[0, 18, 6, 14], [0, 22, 9, 12], [0, 25, 1, 24],
			[0, 27, 11, 16], [0, 23, 7, 26], [1, 19, 7, 13], [1, 23, 10, 15],
			[1, 26, 0, 27], [1, 24, 8, 17], [1, 22, 6, 25], [2, 16, 5, 12],
			[2, 21, 11, 14], [2, 31, 3, 30], [2, 29, 9, 18], [2, 20, 4, 28],
			[3, 17, 4, 15], [3, 20, 8, 13], [3, 28, 2, 29], [3, 30, 10, 19],
			[3, 21, 5, 31], [4, 14, 2, 16], [4, 28, 6, 24], [4, 29, 3, 20],
			[4, 15, 11, 25], [4, 21, 10, 17], [5, 12, 8, 26],
			[5, 20, 9, 16], [5, 13, 3, 17], [5, 31, 7, 27], [5, 30, 2, 21],
			[6, 14, 10, 28], [6, 23, 11, 18], [6, 15, 1, 19],
			[6, 25, 4, 29], [6, 24, 0, 22], [7, 12, 0, 18], [7, 26, 5, 30],
			[7, 27, 1, 23], [7, 13, 9, 31], [7, 22, 8, 19], [8, 13, 1, 22],
			[8, 17, 5, 20], [8, 26, 10, 24], [8, 30, 7, 12], [8, 19, 3, 28],
			[9, 12, 2, 20], [9, 18, 7, 22], [9, 31, 11, 29], [9, 27, 5, 13],
			[9, 16, 0, 25], [10, 15, 3, 21], [10, 19, 6, 23],
			[10, 28, 8, 30], [10, 24, 4, 14], [10, 17, 1, 26],
			[11, 14, 0, 23], [11, 16, 4, 21], [11, 25, 9, 27],
			[11, 29, 6, 15], [11, 18, 2, 31]]
	},
	Polyhedron{
		name:      'SnubCube(dextro}'
		vertexes_: [Vertex{
			x: 0.6212264
			y: -0.3377540
			z: 1.142614
		}, Vertex{
			x: 0.6212264
			y: 0.3377540
			z: -1.142614
		}, Vertex{
			x: -0.6212264
			y: 0.3377540
			z: 1.142614
		}, Vertex{
			x: -0.6212264
			y: -0.3377540
			z: -1.142614
		}, Vertex{
			x: 1.142614
			y: -0.6212264
			z: 0.3377540
		}, Vertex{
			x: 1.142614
			y: 0.6212264
			z: -0.3377540
		}, Vertex{
			x: -1.142614
			y: 0.6212264
			z: 0.3377540
		}, Vertex{
			x: -1.142614
			y: -0.6212264
			z: -0.3377540
		}, Vertex{
			x: 0.3377540
			y: -1.142614
			z: 0.6212264
		}, Vertex{
			x: 0.3377540
			y: 1.142614
			z: -0.6212264
		}, Vertex{
			x: -0.3377540
			y: 1.142614
			z: 0.6212264
		}, Vertex{
			x: -0.3377540
			y: -1.142614
			z: -0.6212264
		}, Vertex{
			x: 0.3377540
			y: 0.6212264
			z: 1.142614
		}, Vertex{
			x: 0.3377540
			y: -0.6212264
			z: -1.142614
		}, Vertex{
			x: -0.3377540
			y: -0.6212264
			z: 1.142614
		}, Vertex{
			x: -0.3377540
			y: 0.6212264
			z: -1.142614
		}, Vertex{
			x: 1.142614
			y: 0.3377540
			z: 0.6212264
		}, Vertex{
			x: 1.142614
			y: -0.3377540
			z: -0.6212264
		}, Vertex{
			x: -1.142614
			y: -0.3377540
			z: 0.6212264
		}, Vertex{
			x: -1.142614
			y: 0.3377540
			z: -0.6212264
		}, Vertex{
			x: 0.6212264
			y: 1.142614
			z: 0.3377540
		}, Vertex{
			x: 0.6212264
			y: -1.142614
			z: -0.3377540
		}, Vertex{
			x: -0.6212264
			y: -1.142614
			z: 0.3377540
		}, Vertex{
			x: -0.6212264
			y: 1.142614
			z: -0.3377540
		}]
		faces:     [[2, 14, 0, 12], [3, 15, 1, 13], [4, 17, 5, 16],
			[7, 18, 6, 19], [8, 22, 11, 21], [9, 23, 10, 20],
			[0, 14, 8], [1, 15, 9], [2, 12, 10], [3, 13, 11],
			[4, 16, 0], [5, 17, 1], [6, 18, 2], [7, 19, 3], [8, 21, 4],
			[9, 20, 5], [10, 23, 6], [11, 22, 7], [12, 0, 16],
			[13, 1, 17], [14, 2, 18], [15, 3, 19], [16, 5, 20],
			[17, 4, 21], [18, 7, 22], [19, 6, 23], [20, 10, 12],
			[21, 11, 13], [22, 8, 14], [23, 9, 15], [8, 4, 0],
			[9, 5, 1], [10, 6, 2], [11, 7, 3], [12, 16, 20], [13, 17, 21],
			[14, 18, 22], [15, 19, 23]]
	},
	Polyhedron{
		name:      'GreatPentagrammicHexecontahedron'
		vertexes_: [Vertex{
			x: -1.438832
			y: 0.5256433
			z: -0.2939417
		}, Vertex{
			x: 1.438832
			y: 0.5256433
			z: 0.2939417
		}, Vertex{
			x: 1.438832
			y: -0.5256433
			z: -0.2939417
		}, Vertex{
			x: -1.438832
			y: -0.5256433
			z: 0.2939417
		}, Vertex{
			x: 0.5256433
			y: -0.2939417
			z: -1.438832
		}, Vertex{
			x: -0.5256433
			y: -0.2939417
			z: 1.438832
		}, Vertex{
			x: -0.5256433
			y: 0.2939417
			z: -1.438832
		}, Vertex{
			x: 0.5256433
			y: 0.2939417
			z: 1.438832
		}, Vertex{
			x: -0.2939417
			y: -1.438832
			z: 0.5256433
		}, Vertex{
			x: 0.2939417
			y: -1.438832
			z: -0.5256433
		}, Vertex{
			x: 0.2939417
			y: 1.438832
			z: 0.5256433
		}, Vertex{
			x: -0.2939417
			y: 1.438832
			z: -0.5256433
		}, Vertex{
			x: 1.457111
			y: 0.0
			z: 0.5565670
		}, Vertex{
			x: 1.457111
			y: 0.0
			z: -0.5565670
		}, Vertex{
			x: -1.457111
			y: 0.0
			z: 0.5565670
		}, Vertex{
			x: -1.457111
			y: 0.0
			z: -0.5565670
		}, Vertex{
			x: 0.0
			y: 0.5565670
			z: 1.457111
		}, Vertex{
			x: 0.0
			y: 0.5565670
			z: -1.457111
		}, Vertex{
			x: 0.0
			y: -0.5565670
			z: 1.457111
		}, Vertex{
			x: 0.0
			y: -0.5565670
			z: -1.457111
		}, Vertex{
			x: 0.5565670
			y: 1.457111
			z: 0.0
		}, Vertex{
			x: -0.5565670
			y: 1.457111
			z: 0.0
		}, Vertex{
			x: 0.5565670
			y: -1.457111
			z: 0.0
		}, Vertex{
			x: -0.5565670
			y: -1.457111
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.3000318
			z: 0.1854299
		}, Vertex{
			x: 0.0
			y: -0.3000318
			z: -0.1854299
		}, Vertex{
			x: 0.0
			y: 0.3000318
			z: 0.1854299
		}, Vertex{
			x: 0.0
			y: 0.3000318
			z: -0.1854299
		}, Vertex{
			x: -0.3000318
			y: 0.1854299
			z: 0.0
		}, Vertex{
			x: 0.3000318
			y: 0.1854299
			z: 0.0
		}, Vertex{
			x: -0.3000318
			y: -0.1854299
			z: 0.0
		}, Vertex{
			x: 0.3000318
			y: -0.1854299
			z: 0.0
		}, Vertex{
			x: 0.1854299
			y: 0.0
			z: -0.3000318
		}, Vertex{
			x: 0.1854299
			y: 0.0
			z: 0.3000318
		}, Vertex{
			x: -0.1854299
			y: 0.0
			z: -0.3000318
		}, Vertex{
			x: -0.1854299
			y: 0.0
			z: 0.3000318
		}, Vertex{
			x: 1.148578
			y: 0.056002
			z: -1.053837
		}, Vertex{
			x: -1.148578
			y: 0.056002
			z: 1.053837
		}, Vertex{
			x: -1.148578
			y: -0.056002
			z: -1.053837
		}, Vertex{
			x: 1.148578
			y: -0.056002
			z: 1.053837
		}, Vertex{
			x: -0.056002
			y: -1.053837
			z: -1.148578
		}, Vertex{
			x: 0.056002
			y: -1.053837
			z: 1.148578
		}, Vertex{
			x: 0.056002
			y: 1.053837
			z: -1.148578
		}, Vertex{
			x: -0.056002
			y: 1.053837
			z: 1.148578
		}, Vertex{
			x: 1.053837
			y: -1.148578
			z: 0.056002
		}, Vertex{
			x: -1.053837
			y: -1.148578
			z: -0.056002
		}, Vertex{
			x: -1.053837
			y: 1.148578
			z: 0.056002
		}, Vertex{
			x: 1.053837
			y: 1.148578
			z: -0.056002
		}, Vertex{
			x: -1.473443
			y: -0.4696413
			z: -0.2033286
		}, Vertex{
			x: 1.473443
			y: -0.4696413
			z: 0.2033286
		}, Vertex{
			x: 1.473443
			y: 0.4696413
			z: -0.2033286
		}, Vertex{
			x: -1.473443
			y: 0.4696413
			z: 0.2033286
		}, Vertex{
			x: -0.4696413
			y: -0.2033286
			z: -1.473443
		}, Vertex{
			x: 0.4696413
			y: -0.2033286
			z: 1.473443
		}, Vertex{
			x: 0.4696413
			y: 0.2033286
			z: -1.473443
		}, Vertex{
			x: -0.4696413
			y: 0.2033286
			z: 1.473443
		}, Vertex{
			x: -0.2033286
			y: -1.473443
			z: -0.4696413
		}, Vertex{
			x: 0.2033286
			y: -1.473443
			z: 0.4696413
		}, Vertex{
			x: 0.2033286
			y: 1.473443
			z: -0.4696413
		}, Vertex{
			x: -0.2033286
			y: 1.473443
			z: 0.4696413
		}, Vertex{
			x: 1.179501
			y: 0.945249
			z: 0.3849946
		}, Vertex{
			x: -1.179501
			y: 0.945249
			z: -0.3849946
		}, Vertex{
			x: -1.179501
			y: -0.945249
			z: 0.3849946
		}, Vertex{
			x: 1.179501
			y: -0.945249
			z: -0.3849946
		}, Vertex{
			x: 0.945249
			y: 0.3849946
			z: 1.179501
		}, Vertex{
			x: -0.945249
			y: 0.3849946
			z: -1.179501
		}, Vertex{
			x: -0.945249
			y: -0.3849946
			z: 1.179501
		}, Vertex{
			x: 0.945249
			y: -0.3849946
			z: -1.179501
		}, Vertex{
			x: 0.3849946
			y: 1.179501
			z: 0.945249
		}, Vertex{
			x: -0.3849946
			y: 1.179501
			z: -0.945249
		}, Vertex{
			x: -0.3849946
			y: -1.179501
			z: 0.945249
		}, Vertex{
			x: 0.3849946
			y: -1.179501
			z: -0.945249
		}, Vertex{
			x: -0.8546358
			y: 0.4196057
			z: 1.235503
		}, Vertex{
			x: 0.8546358
			y: 0.4196057
			z: -1.235503
		}, Vertex{
			x: 0.8546358
			y: -0.4196057
			z: 1.235503
		}, Vertex{
			x: -0.8546358
			y: -0.4196057
			z: -1.235503
		}, Vertex{
			x: -0.4196057
			y: 1.235503
			z: 0.8546358
		}, Vertex{
			x: 0.4196057
			y: 1.235503
			z: -0.8546358
		}, Vertex{
			x: 0.4196057
			y: -1.235503
			z: 0.8546358
		}, Vertex{
			x: -0.4196057
			y: -1.235503
			z: -0.8546358
		}, Vertex{
			x: -1.235503
			y: 0.8546358
			z: 0.4196057
		}, Vertex{
			x: 1.235503
			y: 0.8546358
			z: -0.4196057
		}, Vertex{
			x: 1.235503
			y: -0.8546358
			z: 0.4196057
		}, Vertex{
			x: -1.235503
			y: -0.8546358
			z: -0.4196057
		}, Vertex{
			x: -0.9005442
			y: -0.9005442
			z: -0.9005442
		}, Vertex{
			x: -0.9005442
			y: -0.9005442
			z: 0.9005442
		}, Vertex{
			x: 0.9005442
			y: -0.9005442
			z: -0.9005442
		}, Vertex{
			x: 0.9005442
			y: -0.9005442
			z: 0.9005442
		}, Vertex{
			x: -0.9005442
			y: 0.9005442
			z: -0.9005442
		}, Vertex{
			x: -0.9005442
			y: 0.9005442
			z: 0.9005442
		}, Vertex{
			x: 0.9005442
			y: 0.9005442
			z: -0.9005442
		}, Vertex{
			x: 0.9005442
			y: 0.9005442
			z: 0.9005442
		}]
		faces:     [[24, 0, 2, 14, 36], [24, 36, 72, 86, 76],
			[24, 76, 40, 16, 52], [24, 52, 64, 84, 60], [24, 60, 48, 12, 0],
			[25, 1, 3, 13, 37], [25, 37, 73, 85, 77], [25, 77, 41, 17, 53],
			[25, 53, 65, 87, 61], [25, 61, 49, 15, 1], [26, 2, 0, 12, 38],
			[26, 38, 74, 88, 78], [26, 78, 42, 18, 54], [26, 54, 66, 90, 62],
			[26, 62, 50, 14, 2], [27, 3, 1, 15, 39], [27, 39, 75, 91, 79],
			[27, 79, 43, 19, 55], [27, 55, 67, 89, 63], [27, 63, 51, 13, 3],
			[28, 4, 5, 17, 41], [28, 41, 77, 85, 81], [28, 81, 45, 20, 56],
			[28, 56, 68, 84, 64], [28, 64, 52, 16, 4], [29, 5, 4, 16, 40],
			[29, 40, 76, 86, 80], [29, 80, 44, 21, 57], [29, 57, 69, 87, 65],
			[29, 65, 53, 17, 5], [30, 7, 6, 18, 42], [30, 42, 78, 88, 82],
			[30, 82, 46, 22, 59], [30, 59, 71, 89, 67], [30, 67, 55, 19, 7],
			[31, 6, 7, 19, 43], [31, 43, 79, 91, 83], [31, 83, 47, 23, 58],
			[31, 58, 70, 90, 66], [31, 66, 54, 18, 6], [32, 8, 11, 22, 46],
			[32, 46, 82, 88, 74], [32, 74, 38, 12, 48], [32, 48, 60, 84, 68],
			[32, 68, 56, 20, 8], [33, 11, 8, 20, 45], [33, 45, 81, 85, 73],
			[33, 73, 37, 13, 51], [33, 51, 63, 89, 71], [33, 71, 59, 22, 11],
			[34, 10, 9, 21, 44], [34, 44, 80, 86, 72], [34, 72, 36, 14, 50],
			[34, 50, 62, 90, 70], [34, 70, 58, 23, 10], [35, 9, 10, 23, 47],
			[35, 47, 83, 91, 75], [35, 75, 39, 15, 49], [35, 49, 61, 87, 69],
			[35, 69, 57, 21, 9]]
	},
	Polyhedron{
		name:      'SnubDodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.2015814
			y: -0.2132630
			z: 1.240194
		}, Vertex{
			x: 0.2015814
			y: 0.2132630
			z: -1.240194
		}, Vertex{
			x: -0.2015814
			y: 0.2132630
			z: 1.240194
		}, Vertex{
			x: -0.2015814
			y: -0.2132630
			z: -1.240194
		}, Vertex{
			x: 1.240194
			y: -0.2015814
			z: 0.2132630
		}, Vertex{
			x: 1.240194
			y: 0.2015814
			z: -0.2132630
		}, Vertex{
			x: -1.240194
			y: 0.2015814
			z: 0.2132630
		}, Vertex{
			x: -1.240194
			y: -0.2015814
			z: -0.2132630
		}, Vertex{
			x: 0.2132630
			y: -1.240194
			z: 0.2015814
		}, Vertex{
			x: 0.2132630
			y: 1.240194
			z: -0.2015814
		}, Vertex{
			x: -0.2132630
			y: 1.240194
			z: 0.2015814
		}, Vertex{
			x: -0.2132630
			y: -1.240194
			z: -0.2015814
		}, Vertex{
			x: 0.3114983
			y: 0.3911123
			z: 1.172262
		}, Vertex{
			x: 0.3114983
			y: -0.3911123
			z: -1.172262
		}, Vertex{
			x: -0.3114983
			y: -0.3911123
			z: 1.172262
		}, Vertex{
			x: -0.3114983
			y: 0.3911123
			z: -1.172262
		}, Vertex{
			x: 1.172262
			y: 0.3114983
			z: 0.3911123
		}, Vertex{
			x: 1.172262
			y: -0.3114983
			z: -0.3911123
		}, Vertex{
			x: -1.172262
			y: -0.3114983
			z: 0.3911123
		}, Vertex{
			x: -1.172262
			y: 0.3114983
			z: -0.3911123
		}, Vertex{
			x: 0.3911123
			y: 1.172262
			z: 0.3114983
		}, Vertex{
			x: 0.3911123
			y: -1.172262
			z: -0.3114983
		}, Vertex{
			x: -0.3911123
			y: -1.172262
			z: 0.3114983
		}, Vertex{
			x: -0.3911123
			y: 1.172262
			z: -0.3114983
		}, Vertex{
			x: 0.1099169
			y: -0.7172778
			z: 1.047677
		}, Vertex{
			x: 0.1099169
			y: 0.7172778
			z: -1.047677
		}, Vertex{
			x: -0.1099169
			y: 0.7172778
			z: 1.047677
		}, Vertex{
			x: -0.1099169
			y: -0.7172778
			z: -1.047677
		}, Vertex{
			x: 1.047677
			y: -0.1099169
			z: 0.7172778
		}, Vertex{
			x: 1.047677
			y: 0.1099169
			z: -0.7172778
		}, Vertex{
			x: -1.047677
			y: 0.1099169
			z: 0.7172778
		}, Vertex{
			x: -1.047677
			y: -0.1099169
			z: -0.7172778
		}, Vertex{
			x: 0.7172778
			y: -1.047677
			z: 0.1099169
		}, Vertex{
			x: 0.7172778
			y: 1.047677
			z: -0.1099169
		}, Vertex{
			x: -0.7172778
			y: 1.047677
			z: 0.1099169
		}, Vertex{
			x: -0.7172778
			y: -1.047677
			z: -0.1099169
		}, Vertex{
			x: 0.6565651
			y: -0.5229161
			z: 0.9589985
		}, Vertex{
			x: 0.6565651
			y: 0.5229161
			z: -0.9589985
		}, Vertex{
			x: -0.6565651
			y: 0.5229161
			z: 0.9589985
		}, Vertex{
			x: -0.6565651
			y: -0.5229161
			z: -0.9589985
		}, Vertex{
			x: 0.9589985
			y: -0.6565651
			z: 0.5229161
		}, Vertex{
			x: 0.9589985
			y: 0.6565651
			z: -0.5229161
		}, Vertex{
			x: -0.9589985
			y: 0.6565651
			z: 0.5229161
		}, Vertex{
			x: -0.9589985
			y: -0.6565651
			z: -0.5229161
		}, Vertex{
			x: 0.5229161
			y: -0.9589985
			z: 0.6565651
		}, Vertex{
			x: 0.5229161
			y: 0.9589985
			z: -0.6565651
		}, Vertex{
			x: -0.5229161
			y: 0.9589985
			z: 0.6565651
		}, Vertex{
			x: -0.5229161
			y: -0.9589985
			z: -0.6565651
		}, Vertex{
			x: 0.8344144
			y: 0.4549837
			z: 0.8490816
		}, Vertex{
			x: 0.8344144
			y: -0.4549837
			z: -0.8490816
		}, Vertex{
			x: -0.8344144
			y: -0.4549837
			z: 0.8490816
		}, Vertex{
			x: -0.8344144
			y: 0.4549837
			z: -0.8490816
		}, Vertex{
			x: 0.8490816
			y: 0.8344144
			z: 0.4549837
		}, Vertex{
			x: 0.8490816
			y: -0.8344144
			z: -0.4549837
		}, Vertex{
			x: -0.8490816
			y: -0.8344144
			z: 0.4549837
		}, Vertex{
			x: -0.8490816
			y: 0.8344144
			z: -0.4549837
		}, Vertex{
			x: 0.4549837
			y: 0.8490816
			z: 0.8344144
		}, Vertex{
			x: 0.4549837
			y: -0.8490816
			z: -0.8344144
		}, Vertex{
			x: -0.4549837
			y: -0.8490816
			z: 0.8344144
		}, Vertex{
			x: -0.4549837
			y: 0.8490816
			z: -0.8344144
		}]
		faces:     [[0, 28, 12, 36, 48], [1, 29, 13, 37, 49],
			[2, 30, 14, 38, 50], [3, 31, 15, 39, 51], [4, 32, 17, 40, 53],
			[5, 33, 16, 41, 52], [6, 34, 19, 42, 55], [7, 35, 18, 43, 54],
			[8, 24, 22, 44, 58], [9, 25, 23, 45, 59], [10, 26, 20, 46, 56],
			[11, 27, 21, 47, 57], [0, 26, 42, 18, 58], [1, 27, 43, 19, 59],
			[2, 24, 40, 16, 56], [3, 25, 41, 17, 57], [4, 29, 45, 20, 48],
			[5, 28, 44, 21, 49], [6, 31, 47, 22, 50], [7, 30, 46, 23, 51],
			[8, 35, 39, 13, 53], [9, 34, 38, 12, 52], [10, 33, 37, 15, 55],
			[11, 32, 36, 14, 54], [0, 58, 44], [1, 59, 45], [2, 56, 46],
			[3, 57, 47], [4, 48, 36], [5, 49, 37], [6, 50, 38],
			[7, 51, 39], [8, 53, 40], [9, 52, 41], [10, 55, 42],
			[11, 54, 43], [12, 38, 14], [13, 39, 15], [14, 36, 12],
			[15, 37, 13], [16, 40, 17], [17, 41, 16], [18, 42, 19],
			[19, 43, 18], [20, 45, 23], [21, 44, 22], [22, 47, 21],
			[23, 46, 20], [24, 2, 50], [25, 3, 51], [26, 0, 48],
			[27, 1, 49], [28, 5, 52], [29, 4, 53], [30, 7, 54],
			[31, 6, 55], [32, 11, 57], [33, 10, 56], [34, 9, 59],
			[35, 8, 58], [36, 32, 4], [37, 33, 5], [38, 34, 6],
			[39, 35, 7], [40, 24, 8], [41, 25, 9], [42, 26, 10],
			[43, 27, 11], [44, 28, 0], [45, 29, 1], [46, 30, 2],
			[47, 31, 3], [48, 20, 26], [49, 21, 27], [50, 22, 24],
			[51, 23, 25], [52, 12, 28], [53, 13, 29], [54, 14, 30],
			[55, 15, 31], [56, 16, 33], [57, 17, 32], [58, 18, 35],
			[59, 19, 34]]
	},
	Polyhedron{
		name:      'RhombicDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.060660
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.060660
		}, Vertex{
			x: 1.060660
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.060660
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.060660
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.060660
			z: 0.0
		}, Vertex{
			x: 0.5303301
			y: 0.5303301
			z: 0.5303301
		}, Vertex{
			x: 0.5303301
			y: 0.5303301
			z: -0.5303301
		}, Vertex{
			x: 0.5303301
			y: -0.5303301
			z: 0.5303301
		}, Vertex{
			x: 0.5303301
			y: -0.5303301
			z: -0.5303301
		}, Vertex{
			x: -0.5303301
			y: 0.5303301
			z: 0.5303301
		}, Vertex{
			x: -0.5303301
			y: 0.5303301
			z: -0.5303301
		}, Vertex{
			x: -0.5303301
			y: -0.5303301
			z: 0.5303301
		}, Vertex{
			x: -0.5303301
			y: -0.5303301
			z: -0.5303301
		}]
		faces:     [[6, 0, 8, 2], [6, 2, 7, 4], [6, 4, 10, 0],
			[9, 1, 7, 2], [9, 2, 8, 5], [9, 5, 13, 1], [11, 1, 13, 3],
			[11, 3, 10, 4], [11, 4, 7, 1], [12, 0, 10, 3], [12, 3, 13, 5],
			[12, 5, 8, 0]]
	},
	Polyhedron{
		name:      'DisdyakisDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 2.675417
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -2.675417
		}, Vertex{
			x: 2.675417
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -2.675417
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.675417
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -2.675417
			z: 0.0
		}, Vertex{
			x: 1.640755
			y: 0.0
			z: 1.640755
		}, Vertex{
			x: 1.640755
			y: 0.0
			z: -1.640755
		}, Vertex{
			x: -1.640755
			y: 0.0
			z: 1.640755
		}, Vertex{
			x: -1.640755
			y: 0.0
			z: -1.640755
		}, Vertex{
			x: 1.640755
			y: 1.640755
			z: 0.0
		}, Vertex{
			x: 1.640755
			y: -1.640755
			z: 0.0
		}, Vertex{
			x: -1.640755
			y: 1.640755
			z: 0.0
		}, Vertex{
			x: -1.640755
			y: -1.640755
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.640755
			z: 1.640755
		}, Vertex{
			x: 0.0
			y: 1.640755
			z: -1.640755
		}, Vertex{
			x: 0.0
			y: -1.640755
			z: 1.640755
		}, Vertex{
			x: 0.0
			y: -1.640755
			z: -1.640755
		}, Vertex{
			x: 1.414214
			y: 1.414214
			z: 1.414214
		}, Vertex{
			x: 1.414214
			y: 1.414214
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: -1.414214
			z: 1.414214
		}, Vertex{
			x: 1.414214
			y: -1.414214
			z: -1.414214
		}, Vertex{
			x: -1.414214
			y: 1.414214
			z: 1.414214
		}, Vertex{
			x: -1.414214
			y: 1.414214
			z: -1.414214
		}, Vertex{
			x: -1.414214
			y: -1.414214
			z: 1.414214
		}, Vertex{
			x: -1.414214
			y: -1.414214
			z: -1.414214
		}]
		faces:     [[0, 6, 18], [0, 18, 14], [0, 14, 22], [0, 22, 8],
			[0, 8, 24], [0, 24, 16], [0, 16, 20], [0, 20, 6],
			[1, 7, 21], [1, 21, 17], [1, 17, 25], [1, 25, 9],
			[1, 9, 23], [1, 23, 15], [1, 15, 19], [1, 19, 7],
			[2, 6, 20], [2, 20, 11], [2, 11, 21], [2, 21, 7],
			[2, 7, 19], [2, 19, 10], [2, 10, 18], [2, 18, 6],
			[3, 8, 22], [3, 22, 12], [3, 12, 23], [3, 23, 9],
			[3, 9, 25], [3, 25, 13], [3, 13, 24], [3, 24, 8],
			[4, 10, 19], [4, 19, 15], [4, 15, 23], [4, 23, 12],
			[4, 12, 22], [4, 22, 14], [4, 14, 18], [4, 18, 10],
			[5, 11, 20], [5, 20, 16], [5, 16, 24], [5, 24, 13],
			[5, 13, 25], [5, 25, 17], [5, 17, 21], [5, 21, 11]]
	},
	Polyhedron{
		name:      'SmallIcosihemidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: -1.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: -1.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: -1.309017
			z: -0.5
		}]
		faces:     [[0, 6, 22, 23, 7, 1, 13, 29, 28, 12], [0, 8, 24, 25, 9, 1, 11, 27, 26, 10],
			[2, 14, 6, 10, 18, 3, 21, 13, 9, 17], [2, 15, 7, 11, 19, 3, 20, 12, 8, 16],
			[4, 22, 14, 16, 24, 5, 29, 21, 19, 27], [4, 23, 15, 17, 25, 5, 28, 20, 18, 26],
			[0, 6, 10], [0, 12, 8], [1, 9, 13], [1, 11, 7], [14, 16, 2],
			[14, 22, 6], [17, 15, 2], [17, 25, 9], [19, 21, 3],
			[19, 27, 11], [20, 18, 3], [20, 28, 12], [23, 4, 22],
			[23, 15, 7], [24, 5, 25], [24, 16, 8], [26, 4, 27],
			[26, 18, 10], [29, 5, 28], [29, 21, 13]]
	},
	Polyhedron{
		name:      'Rhombicosacron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.341641
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.341641
		}, Vertex{
			x: 1.341641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.341641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.341641
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.341641
			z: 0.0
		}, Vertex{
			x: 0.4145898
			y: 0.6708204
			z: 1.085410
		}, Vertex{
			x: 0.4145898
			y: 0.6708204
			z: -1.085410
		}, Vertex{
			x: 0.4145898
			y: -0.6708204
			z: 1.085410
		}, Vertex{
			x: 0.4145898
			y: -0.6708204
			z: -1.085410
		}, Vertex{
			x: -0.4145898
			y: 0.6708204
			z: 1.085410
		}, Vertex{
			x: -0.4145898
			y: 0.6708204
			z: -1.085410
		}, Vertex{
			x: -0.4145898
			y: -0.6708204
			z: 1.085410
		}, Vertex{
			x: -0.4145898
			y: -0.6708204
			z: -1.085410
		}, Vertex{
			x: 1.085410
			y: 0.4145898
			z: 0.6708204
		}, Vertex{
			x: 1.085410
			y: 0.4145898
			z: -0.6708204
		}, Vertex{
			x: 1.085410
			y: -0.4145898
			z: 0.6708204
		}, Vertex{
			x: 1.085410
			y: -0.4145898
			z: -0.6708204
		}, Vertex{
			x: -1.085410
			y: 0.4145898
			z: 0.6708204
		}, Vertex{
			x: -1.085410
			y: 0.4145898
			z: -0.6708204
		}, Vertex{
			x: -1.085410
			y: -0.4145898
			z: 0.6708204
		}, Vertex{
			x: -1.085410
			y: -0.4145898
			z: -0.6708204
		}, Vertex{
			x: 0.6708204
			y: 1.085410
			z: 0.4145898
		}, Vertex{
			x: 0.6708204
			y: 1.085410
			z: -0.4145898
		}, Vertex{
			x: 0.6708204
			y: -1.085410
			z: 0.4145898
		}, Vertex{
			x: 0.6708204
			y: -1.085410
			z: -0.4145898
		}, Vertex{
			x: -0.6708204
			y: 1.085410
			z: 0.4145898
		}, Vertex{
			x: -0.6708204
			y: 1.085410
			z: -0.4145898
		}, Vertex{
			x: -0.6708204
			y: -1.085410
			z: 0.4145898
		}, Vertex{
			x: -0.6708204
			y: -1.085410
			z: -0.4145898
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[0, 16, 8, 22], [0, 28, 44, 18], [0, 32, 6, 12],
			[1, 16, 10, 19], [1, 33, 49, 23], [1, 29, 5, 13],
			[2, 17, 11, 20], [2, 30, 46, 24], [2, 26, 4, 12],
			[3, 17, 9, 25], [3, 27, 43, 21], [3, 31, 7, 13], [4, 12, 0, 28],
			[4, 35, 43, 26], [4, 37, 9, 14], [5, 13, 3, 27], [5, 36, 44, 29],
			[5, 34, 8, 14], [6, 12, 2, 30], [6, 41, 49, 32], [6, 39, 10, 15],
			[7, 13, 1, 33], [7, 38, 46, 31], [7, 40, 11, 15],
			[8, 14, 4, 35], [8, 22, 46, 34], [8, 23, 1, 16], [9, 14, 5, 36],
			[9, 25, 49, 37], [9, 24, 2, 17], [10, 15, 7, 38],
			[10, 19, 43, 39], [10, 18, 0, 16], [11, 15, 6, 41],
			[11, 20, 44, 40], [11, 21, 3, 17], [42, 20, 2, 26],
			[42, 38, 10, 18], [42, 27, 5, 34], [43, 21, 45, 19],
			[43, 26, 42, 27], [43, 39, 47, 35], [44, 18, 42, 20],
			[44, 29, 45, 28], [44, 40, 48, 36], [45, 19, 1, 29],
			[45, 41, 11, 21], [45, 28, 4, 37], [46, 24, 48, 22],
			[46, 31, 47, 30], [46, 34, 42, 38], [47, 25, 3, 31],
			[47, 35, 8, 23], [47, 30, 6, 39], [48, 22, 0, 32],
			[48, 36, 9, 24], [48, 33, 7, 40], [49, 23, 47, 25],
			[49, 32, 48, 33], [49, 37, 45, 41]]
	},
	Polyhedron{
		name:      'Cube'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.5
		}]
		faces:     [[0, 1, 5, 4], [0, 4, 6, 2], [0, 2, 3, 1],
			[7, 3, 2, 6], [7, 6, 4, 5], [7, 5, 1, 3]]
	},
	Polyhedron{
		name:      'GreatDeltoidalIcositetrahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.414214
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: -0.3693981
			y: -0.3693981
			z: -0.3693981
		}, Vertex{
			x: -0.3693981
			y: -0.3693981
			z: 0.3693981
		}, Vertex{
			x: -0.3693981
			y: 0.3693981
			z: -0.3693981
		}, Vertex{
			x: -0.3693981
			y: 0.3693981
			z: 0.3693981
		}, Vertex{
			x: 0.3693981
			y: -0.3693981
			z: -0.3693981
		}, Vertex{
			x: 0.3693981
			y: -0.3693981
			z: 0.3693981
		}, Vertex{
			x: 0.3693981
			y: 0.3693981
			z: -0.3693981
		}, Vertex{
			x: 0.3693981
			y: 0.3693981
			z: 0.3693981
		}]
		faces:     [[0, 6, 18, 14], [0, 14, 22, 8], [0, 8, 24, 16],
			[0, 16, 20, 6], [1, 9, 23, 15], [1, 15, 19, 7], [1, 7, 21, 17],
			[1, 17, 25, 9], [2, 7, 19, 10], [2, 10, 18, 6], [2, 6, 20, 11],
			[2, 11, 21, 7], [3, 8, 22, 12], [3, 12, 23, 9], [3, 9, 25, 13],
			[3, 13, 24, 8], [4, 10, 19, 15], [4, 15, 23, 12],
			[4, 12, 22, 14], [4, 14, 18, 10], [5, 11, 20, 16],
			[5, 16, 24, 13], [5, 13, 25, 17], [5, 17, 21, 11]]
	},
	Polyhedron{
		name:      'SnubIcosidodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.1053988
			y: -0.1849619
			z: 1.106607
		}, Vertex{
			x: 0.1053988
			y: 0.1849619
			z: -1.106607
		}, Vertex{
			x: -0.1053988
			y: 0.1849619
			z: 1.106607
		}, Vertex{
			x: -0.1053988
			y: -0.1849619
			z: -1.106607
		}, Vertex{
			x: 1.106607
			y: -0.1053988
			z: 0.1849619
		}, Vertex{
			x: 1.106607
			y: 0.1053988
			z: -0.1849619
		}, Vertex{
			x: -1.106607
			y: 0.1053988
			z: 0.1849619
		}, Vertex{
			x: -1.106607
			y: -0.1053988
			z: -0.1849619
		}, Vertex{
			x: 0.1849619
			y: -1.106607
			z: 0.1053988
		}, Vertex{
			x: 0.1849619
			y: 1.106607
			z: -0.1053988
		}, Vertex{
			x: -0.1849619
			y: 1.106607
			z: 0.1053988
		}, Vertex{
			x: -0.1849619
			y: -1.106607
			z: -0.1053988
		}, Vertex{
			x: 0.2450224
			y: 0.4108777
			z: 1.020315
		}, Vertex{
			x: 0.2450224
			y: -0.4108777
			z: -1.020315
		}, Vertex{
			x: -0.2450224
			y: -0.4108777
			z: 1.020315
		}, Vertex{
			x: -0.2450224
			y: 0.4108777
			z: -1.020315
		}, Vertex{
			x: 1.020315
			y: 0.2450224
			z: 0.4108777
		}, Vertex{
			x: 1.020315
			y: -0.2450224
			z: -0.4108777
		}, Vertex{
			x: -1.020315
			y: -0.2450224
			z: 0.4108777
		}, Vertex{
			x: -1.020315
			y: 0.2450224
			z: -0.4108777
		}, Vertex{
			x: 0.4108777
			y: 1.020315
			z: 0.2450224
		}, Vertex{
			x: 0.4108777
			y: -1.020315
			z: -0.2450224
		}, Vertex{
			x: -0.4108777
			y: -1.020315
			z: 0.2450224
		}, Vertex{
			x: -0.4108777
			y: 1.020315
			z: -0.2450224
		}, Vertex{
			x: 0.1396236
			y: -0.5814166
			z: 0.9551749
		}, Vertex{
			x: 0.1396236
			y: 0.5814166
			z: -0.9551749
		}, Vertex{
			x: -0.1396236
			y: 0.5814166
			z: 0.9551749
		}, Vertex{
			x: -0.1396236
			y: -0.5814166
			z: -0.9551749
		}, Vertex{
			x: 0.9551749
			y: -0.1396236
			z: 0.5814166
		}, Vertex{
			x: 0.9551749
			y: 0.1396236
			z: -0.5814166
		}, Vertex{
			x: -0.9551749
			y: 0.1396236
			z: 0.5814166
		}, Vertex{
			x: -0.9551749
			y: -0.1396236
			z: -0.5814166
		}, Vertex{
			x: 0.5814166
			y: -0.9551749
			z: 0.1396236
		}, Vertex{
			x: 0.5814166
			y: 0.9551749
			z: -0.1396236
		}, Vertex{
			x: -0.5814166
			y: 0.9551749
			z: 0.1396236
		}, Vertex{
			x: -0.5814166
			y: -0.9551749
			z: -0.1396236
		}, Vertex{
			x: 0.5442971
			y: -0.5251905
			z: 0.8353529
		}, Vertex{
			x: 0.5442971
			y: 0.5251905
			z: -0.8353529
		}, Vertex{
			x: -0.5442971
			y: 0.5251905
			z: 0.8353529
		}, Vertex{
			x: -0.5442971
			y: -0.5251905
			z: -0.8353529
		}, Vertex{
			x: 0.8353529
			y: -0.5442971
			z: 0.5251905
		}, Vertex{
			x: 0.8353529
			y: 0.5442971
			z: -0.5251905
		}, Vertex{
			x: -0.8353529
			y: 0.5442971
			z: 0.5251905
		}, Vertex{
			x: -0.8353529
			y: -0.5442971
			z: -0.5251905
		}, Vertex{
			x: 0.5251905
			y: -0.8353529
			z: 0.5442971
		}, Vertex{
			x: 0.5251905
			y: 0.8353529
			z: -0.5442971
		}, Vertex{
			x: -0.5251905
			y: 0.8353529
			z: 0.5442971
		}, Vertex{
			x: -0.5251905
			y: -0.8353529
			z: -0.5442971
		}, Vertex{
			x: 0.4388984
			y: 0.6957293
			z: 0.7702129
		}, Vertex{
			x: 0.4388984
			y: -0.6957293
			z: -0.7702129
		}, Vertex{
			x: -0.4388984
			y: -0.6957293
			z: 0.7702129
		}, Vertex{
			x: -0.4388984
			y: 0.6957293
			z: -0.7702129
		}, Vertex{
			x: 0.7702129
			y: 0.4388984
			z: 0.6957293
		}, Vertex{
			x: 0.7702129
			y: -0.4388984
			z: -0.6957293
		}, Vertex{
			x: -0.7702129
			y: -0.4388984
			z: 0.6957293
		}, Vertex{
			x: -0.7702129
			y: 0.4388984
			z: -0.6957293
		}, Vertex{
			x: 0.6957293
			y: 0.7702129
			z: 0.4388984
		}, Vertex{
			x: 0.6957293
			y: -0.7702129
			z: -0.4388984
		}, Vertex{
			x: -0.6957293
			y: -0.7702129
			z: 0.4388984
		}, Vertex{
			x: -0.6957293
			y: 0.7702129
			z: -0.4388984
		}]
		faces:     [[0, 52, 36, 12, 28], [1, 53, 37, 13, 29],
			[2, 54, 38, 14, 30], [3, 55, 39, 15, 31], [4, 57, 40, 17, 32],
			[5, 56, 41, 16, 33], [6, 59, 42, 19, 34], [7, 58, 43, 18, 35],
			[8, 50, 44, 22, 24], [9, 51, 45, 23, 25], [10, 48, 46, 20, 26],
			[11, 49, 47, 21, 27], [0, 54, 35, 21, 40], [1, 55, 34, 20, 41],
			[2, 52, 33, 23, 42], [3, 53, 32, 22, 43], [4, 56, 26, 14, 44],
			[5, 57, 27, 15, 45], [6, 58, 24, 12, 46], [7, 59, 25, 13, 47],
			[8, 49, 29, 16, 36], [9, 48, 28, 17, 37], [10, 51, 31, 18, 38],
			[11, 50, 30, 19, 39], [0, 28, 48], [1, 29, 49], [2, 30, 50],
			[3, 31, 51], [4, 32, 53], [5, 33, 52], [6, 34, 55],
			[7, 35, 54], [8, 24, 58], [9, 25, 59], [10, 26, 56],
			[11, 27, 57], [12, 20, 46], [13, 21, 47], [14, 22, 44],
			[15, 23, 45], [16, 12, 36], [17, 13, 37], [18, 14, 38],
			[19, 15, 39], [20, 16, 41], [21, 17, 40], [22, 18, 43],
			[23, 19, 42], [24, 28, 12], [25, 29, 13], [26, 30, 14],
			[27, 31, 15], [28, 32, 17], [29, 33, 16], [30, 34, 19],
			[31, 35, 18], [32, 24, 22], [33, 25, 23], [34, 26, 20],
			[35, 27, 21], [36, 50, 8], [37, 51, 9], [38, 48, 10],
			[39, 49, 11], [40, 52, 0], [41, 53, 1], [42, 54, 2],
			[43, 55, 3], [44, 57, 4], [45, 56, 5], [46, 59, 6],
			[47, 58, 7], [48, 9, 46], [49, 8, 47], [50, 11, 44],
			[51, 10, 45], [52, 2, 36], [53, 3, 37], [54, 0, 38],
			[55, 1, 39], [56, 4, 41], [57, 5, 40], [58, 6, 43],
			[59, 7, 42], [0, 48, 38], [1, 49, 39], [2, 50, 36],
			[3, 51, 37], [4, 53, 41], [5, 52, 40], [6, 55, 43],
			[7, 54, 42], [8, 58, 47], [9, 59, 46], [10, 56, 45],
			[11, 57, 44], [12, 16, 20], [13, 17, 21], [14, 18, 22],
			[15, 19, 23], [24, 32, 28], [25, 33, 29], [26, 34, 30],
			[27, 35, 31]]
	},
	Polyhedron{
		name:      'GreatDeltoidalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: -2.236068
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 2.236068
		}, Vertex{
			x: 0.0
			y: -2.236068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.236068
			z: 0.0
		}, Vertex{
			x: -2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.5801787
			y: 0.0
			z: 0.2216086
		}, Vertex{
			x: 0.5801787
			y: 0.0
			z: -0.2216086
		}, Vertex{
			x: -0.5801787
			y: 0.0
			z: 0.2216086
		}, Vertex{
			x: -0.5801787
			y: 0.0
			z: -0.2216086
		}, Vertex{
			x: 0.0
			y: 0.2216086
			z: 0.5801787
		}, Vertex{
			x: 0.0
			y: 0.2216086
			z: -0.5801787
		}, Vertex{
			x: 0.0
			y: -0.2216086
			z: 0.5801787
		}, Vertex{
			x: 0.0
			y: -0.2216086
			z: -0.5801787
		}, Vertex{
			x: 0.2216086
			y: 0.5801787
			z: 0.0
		}, Vertex{
			x: -0.2216086
			y: 0.5801787
			z: 0.0
		}, Vertex{
			x: 0.2216086
			y: -0.5801787
			z: 0.0
		}, Vertex{
			x: -0.2216086
			y: -0.5801787
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.4606553
			z: -0.2847007
		}, Vertex{
			x: 0.0
			y: 0.4606553
			z: 0.2847007
		}, Vertex{
			x: 0.0
			y: -0.4606553
			z: -0.2847007
		}, Vertex{
			x: 0.0
			y: -0.4606553
			z: 0.2847007
		}, Vertex{
			x: 0.4606553
			y: -0.2847007
			z: 0.0
		}, Vertex{
			x: -0.4606553
			y: -0.2847007
			z: 0.0
		}, Vertex{
			x: 0.4606553
			y: 0.2847007
			z: 0.0
		}, Vertex{
			x: -0.4606553
			y: 0.2847007
			z: 0.0
		}, Vertex{
			x: -0.2847007
			y: 0.0
			z: 0.4606553
		}, Vertex{
			x: -0.2847007
			y: 0.0
			z: -0.4606553
		}, Vertex{
			x: 0.2847007
			y: 0.0
			z: 0.4606553
		}, Vertex{
			x: 0.2847007
			y: 0.0
			z: -0.4606553
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: -0.3585702
			y: -0.3585702
			z: -0.3585702
		}, Vertex{
			x: -0.3585702
			y: -0.3585702
			z: 0.3585702
		}, Vertex{
			x: 0.3585702
			y: -0.3585702
			z: -0.3585702
		}, Vertex{
			x: 0.3585702
			y: -0.3585702
			z: 0.3585702
		}, Vertex{
			x: -0.3585702
			y: 0.3585702
			z: -0.3585702
		}, Vertex{
			x: -0.3585702
			y: 0.3585702
			z: 0.3585702
		}, Vertex{
			x: 0.3585702
			y: 0.3585702
			z: -0.3585702
		}, Vertex{
			x: 0.3585702
			y: 0.3585702
			z: 0.3585702
		}]
		faces:     [[18, 0, 8, 32], [18, 32, 56, 40], [18, 40, 10, 38],
			[18, 38, 54, 30], [18, 30, 6, 0], [19, 1, 7, 31],
			[19, 31, 55, 39], [19, 39, 11, 41], [19, 41, 57, 33],
			[19, 33, 9, 1], [20, 0, 6, 34], [20, 34, 58, 42],
			[20, 42, 12, 44], [20, 44, 60, 36], [20, 36, 8, 0],
			[21, 1, 9, 37], [21, 37, 61, 45], [21, 45, 13, 43],
			[21, 43, 59, 35], [21, 35, 7, 1], [22, 2, 11, 39],
			[22, 39, 55, 47], [22, 47, 14, 46], [22, 46, 54, 38],
			[22, 38, 10, 2], [23, 2, 10, 40], [23, 40, 56, 48],
			[23, 48, 15, 49], [23, 49, 57, 41], [23, 41, 11, 2],
			[24, 3, 12, 42], [24, 42, 58, 50], [24, 50, 16, 51],
			[24, 51, 59, 43], [24, 43, 13, 3], [25, 3, 13, 45],
			[25, 45, 61, 53], [25, 53, 17, 52], [25, 52, 60, 44],
			[25, 44, 12, 3], [26, 4, 16, 50], [26, 50, 58, 34],
			[26, 34, 6, 30], [26, 30, 54, 46], [26, 46, 14, 4],
			[27, 4, 14, 47], [27, 47, 55, 31], [27, 31, 7, 35],
			[27, 35, 59, 51], [27, 51, 16, 4], [28, 5, 15, 48],
			[28, 48, 56, 32], [28, 32, 8, 36], [28, 36, 60, 52],
			[28, 52, 17, 5], [29, 5, 17, 53], [29, 53, 61, 37],
			[29, 37, 9, 33], [29, 33, 57, 49], [29, 49, 15, 5]]
	},
	Polyhedron{
		name:      'Tetrahedron'
		vertexes_: [Vertex{
			x: 0.3535534
			y: -0.3535534
			z: 0.3535534
		}, Vertex{
			x: 0.3535534
			y: 0.3535534
			z: -0.3535534
		}, Vertex{
			x: -0.3535534
			y: 0.3535534
			z: 0.3535534
		}, Vertex{
			x: -0.3535534
			y: -0.3535534
			z: -0.3535534
		}]
		faces:     [[0, 1, 2], [1, 0, 3], [2, 3, 0], [3, 2, 1]]
	},
	Polyhedron{
		name:      'SmallDodecahemidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: -1.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: -1.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: -1.309017
			z: -0.5
		}]
		faces:     [[0, 6, 22, 23, 7, 1, 13, 29, 28, 12], [0, 8, 24, 25, 9, 1, 11, 27, 26, 10],
			[2, 14, 6, 10, 18, 3, 21, 13, 9, 17], [2, 15, 7, 11, 19, 3, 20, 12, 8, 16],
			[4, 22, 14, 16, 24, 5, 29, 21, 19, 27], [4, 23, 15, 17, 25, 5, 28, 20, 18, 26],
			[0, 8, 16, 14, 6], [0, 10, 18, 20, 12], [1, 7, 15, 17, 9],
			[1, 13, 21, 19, 11], [2, 15, 23, 22, 14], [2, 16, 24, 25, 17],
			[3, 18, 26, 27, 19], [3, 21, 29, 28, 20], [4, 23, 7, 11, 27],
			[4, 26, 10, 6, 22], [5, 24, 8, 12, 28], [5, 29, 13, 9, 25]]
	},
	Polyhedron{
		name:      'GreatDodecicosahedron'
		vertexes_: [Vertex{
			x: -0.809017
			y: 0.5
			z: -0.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: 0.618034
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: -0.618034
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: 0.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: -0.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: 0.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: -0.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: 0.618034
		}, Vertex{
			x: 0.5
			y: -0.618034
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: -0.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: -0.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: -0.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: 0.618034
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: 0.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: 0.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: 0.618034
			z: 0.809017
		}, Vertex{
			x: -0.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: -0.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: 0.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: 0.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: -0.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: 0.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: 0.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: -1.118034
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: 1.118034
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: 1.118034
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: -1.118034
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: 1.118034
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: -1.118034
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: 1.118034
		}, Vertex{
			x: 0.1909830
			y: -1.118034
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: -1.118034
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: 1.118034
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: 1.118034
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 1.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: 1.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: 1.0
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: 1.0
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: -1.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: -1.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: -1.0
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: -1.0
			z: -0.1909830
		}, Vertex{
			x: 1.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: 1.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: -1.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: -1.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: 1.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: 1.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: -1.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: -1.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: 1.0
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: -1.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: 1.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: -1.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: 1.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: -1.0
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: 1.0
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: -1.0
		}]
		faces:     [[0, 4, 30, 14, 51, 59, 55, 47, 10, 28], [0, 38, 46, 47, 39, 1, 25, 21, 20, 24],
			[2, 26, 22, 23, 27, 3, 37, 45, 44, 36], [2, 28, 8, 45, 53, 57, 49, 12, 30, 6],
			[5, 1, 29, 11, 46, 54, 58, 50, 15, 31], [5, 43, 51, 50, 42, 4, 24, 16, 17, 25],
			[7, 27, 19, 18, 26, 6, 40, 48, 49, 41], [7, 31, 13, 48, 56, 52, 44, 9, 29, 3],
			[33, 11, 9, 32, 16, 56, 40, 42, 58, 18], [33, 19, 59, 43, 41, 57, 17, 32, 8, 10],
			[34, 13, 15, 35, 22, 54, 38, 36, 52, 20], [34, 21, 53, 37, 39, 55, 23, 35, 14, 12],
			[0, 4, 42, 58, 54, 38], [0, 28, 8, 32, 16, 24], [3, 7, 41, 57, 53, 37],
			[3, 29, 11, 33, 19, 27], [17, 32, 9, 29, 1, 25], [17, 57, 49, 48, 56, 16],
			[18, 33, 10, 28, 2, 26], [18, 58, 50, 51, 59, 19],
			[34, 12, 30, 4, 24, 20], [34, 21, 25, 5, 31, 13],
			[35, 15, 31, 7, 27, 23], [35, 22, 26, 6, 30, 14],
			[40, 6, 2, 36, 52, 56], [40, 48, 13, 15, 50, 42],
			[43, 5, 1, 39, 55, 59], [43, 51, 14, 12, 49, 41],
			[44, 36, 38, 46, 11, 9], [44, 45, 53, 21, 20, 52],
			[47, 39, 37, 45, 8, 10], [47, 46, 54, 22, 23, 55]]
	},
	Polyhedron{
		name:      'GreatRetrosnubIcosidodecahedron'
		vertexes_: [Vertex{
			x: -0.1715724
			y: 0.4696413
			z: 0.2939417
		}, Vertex{
			x: 0.1715724
			y: 0.4696413
			z: -0.2939417
		}, Vertex{
			x: 0.1715724
			y: -0.4696413
			z: 0.2939417
		}, Vertex{
			x: -0.1715724
			y: -0.4696413
			z: -0.2939417
		}, Vertex{
			x: 0.4696413
			y: 0.2939417
			z: -0.1715724
		}, Vertex{
			x: -0.4696413
			y: 0.2939417
			z: 0.1715724
		}, Vertex{
			x: -0.4696413
			y: -0.2939417
			z: -0.1715724
		}, Vertex{
			x: 0.4696413
			y: -0.2939417
			z: 0.1715724
		}, Vertex{
			x: 0.2939417
			y: -0.1715724
			z: 0.4696413
		}, Vertex{
			x: -0.2939417
			y: -0.1715724
			z: -0.4696413
		}, Vertex{
			x: -0.2939417
			y: 0.1715724
			z: 0.4696413
		}, Vertex{
			x: 0.2939417
			y: 0.1715724
			z: -0.4696413
		}, Vertex{
			x: -0.1532930
			y: -0.056002
			z: -0.5565670
		}, Vertex{
			x: 0.1532930
			y: -0.056002
			z: 0.5565670
		}, Vertex{
			x: 0.1532930
			y: 0.056002
			z: -0.5565670
		}, Vertex{
			x: -0.1532930
			y: 0.056002
			z: 0.5565670
		}, Vertex{
			x: 0.056002
			y: -0.5565670
			z: 0.1532930
		}, Vertex{
			x: -0.056002
			y: -0.5565670
			z: -0.1532930
		}, Vertex{
			x: -0.056002
			y: 0.5565670
			z: 0.1532930
		}, Vertex{
			x: 0.056002
			y: 0.5565670
			z: -0.1532930
		}, Vertex{
			x: 0.5565670
			y: 0.1532930
			z: -0.056002
		}, Vertex{
			x: -0.5565670
			y: 0.1532930
			z: 0.056002
		}, Vertex{
			x: -0.5565670
			y: -0.1532930
			z: -0.056002
		}, Vertex{
			x: 0.5565670
			y: -0.1532930
			z: 0.056002
		}, Vertex{
			x: -0.1369612
			y: -0.5256433
			z: 0.2033286
		}, Vertex{
			x: 0.1369612
			y: -0.5256433
			z: -0.2033286
		}, Vertex{
			x: 0.1369612
			y: 0.5256433
			z: 0.2033286
		}, Vertex{
			x: -0.1369612
			y: 0.5256433
			z: -0.2033286
		}, Vertex{
			x: -0.5256433
			y: 0.2033286
			z: -0.1369612
		}, Vertex{
			x: 0.5256433
			y: 0.2033286
			z: 0.1369612
		}, Vertex{
			x: 0.5256433
			y: -0.2033286
			z: -0.1369612
		}, Vertex{
			x: -0.5256433
			y: -0.2033286
			z: 0.1369612
		}, Vertex{
			x: 0.2033286
			y: -0.1369612
			z: -0.5256433
		}, Vertex{
			x: -0.2033286
			y: -0.1369612
			z: 0.5256433
		}, Vertex{
			x: -0.2033286
			y: 0.1369612
			z: -0.5256433
		}, Vertex{
			x: 0.2033286
			y: 0.1369612
			z: 0.5256433
		}, Vertex{
			x: 0.4309030
			y: 0.05003555
			z: -0.3849946
		}, Vertex{
			x: -0.4309030
			y: 0.05003555
			z: 0.3849946
		}, Vertex{
			x: -0.4309030
			y: -0.05003555
			z: -0.3849946
		}, Vertex{
			x: 0.4309030
			y: -0.05003555
			z: 0.3849946
		}, Vertex{
			x: 0.05003555
			y: -0.3849946
			z: 0.4309030
		}, Vertex{
			x: -0.05003555
			y: -0.3849946
			z: -0.4309030
		}, Vertex{
			x: -0.05003555
			y: 0.3849946
			z: 0.4309030
		}, Vertex{
			x: 0.05003555
			y: 0.3849946
			z: -0.4309030
		}, Vertex{
			x: -0.3849946
			y: 0.4309030
			z: 0.05003555
		}, Vertex{
			x: 0.3849946
			y: 0.4309030
			z: -0.05003555
		}, Vertex{
			x: 0.3849946
			y: -0.4309030
			z: 0.05003555
		}, Vertex{
			x: -0.3849946
			y: -0.4309030
			z: -0.05003555
		}, Vertex{
			x: 0.4196057
			y: 0.3749010
			z: 0.1406487
		}, Vertex{
			x: -0.4196057
			y: 0.3749010
			z: -0.1406487
		}, Vertex{
			x: -0.4196057
			y: -0.3749010
			z: 0.1406487
		}, Vertex{
			x: 0.4196057
			y: -0.3749010
			z: -0.1406487
		}, Vertex{
			x: -0.3749010
			y: 0.1406487
			z: -0.4196057
		}, Vertex{
			x: 0.3749010
			y: 0.1406487
			z: 0.4196057
		}, Vertex{
			x: 0.3749010
			y: -0.1406487
			z: -0.4196057
		}, Vertex{
			x: -0.3749010
			y: -0.1406487
			z: 0.4196057
		}, Vertex{
			x: -0.1406487
			y: -0.4196057
			z: 0.3749010
		}, Vertex{
			x: 0.1406487
			y: -0.4196057
			z: -0.3749010
		}, Vertex{
			x: 0.1406487
			y: 0.4196057
			z: 0.3749010
		}, Vertex{
			x: -0.1406487
			y: 0.4196057
			z: -0.3749010
		}]
		faces:     [[0, 36, 28, 48, 12], [1, 37, 29, 49, 13],
			[2, 38, 30, 50, 14], [3, 39, 31, 51, 15], [4, 40, 32, 53, 17],
			[5, 41, 33, 52, 16], [6, 42, 34, 55, 19], [7, 43, 35, 54, 18],
			[8, 44, 24, 58, 22], [9, 45, 25, 59, 23], [10, 46, 26, 56, 20],
			[11, 47, 27, 57, 21], [0, 2, 14], [1, 3, 15], [2, 0, 12],
			[3, 1, 13], [4, 5, 16], [5, 4, 17], [6, 7, 18], [7, 6, 19],
			[8, 11, 21], [9, 10, 20], [10, 9, 23], [11, 8, 22],
			[12, 48, 56], [13, 49, 57], [14, 50, 58], [15, 51, 59],
			[16, 52, 48], [17, 53, 49], [18, 54, 50], [19, 55, 51],
			[20, 56, 52], [21, 57, 53], [22, 58, 54], [23, 59, 55],
			[24, 44, 36], [25, 45, 37], [26, 46, 38], [27, 47, 39],
			[28, 36, 40], [29, 37, 41], [30, 38, 42], [31, 39, 43],
			[32, 40, 44], [33, 41, 45], [34, 42, 46], [35, 43, 47],
			[36, 0, 24], [37, 1, 25], [38, 2, 26], [39, 3, 27],
			[40, 4, 28], [41, 5, 29], [42, 6, 30], [43, 7, 31],
			[44, 8, 32], [45, 9, 33], [46, 10, 34], [47, 11, 35],
			[48, 28, 16], [49, 29, 17], [50, 30, 18], [51, 31, 19],
			[52, 33, 20], [53, 32, 21], [54, 35, 22], [55, 34, 23],
			[56, 26, 12], [57, 27, 13], [58, 24, 14], [59, 25, 15],
			[24, 0, 14], [25, 1, 15], [26, 2, 12], [27, 3, 13],
			[28, 4, 16], [29, 5, 17], [30, 6, 18], [31, 7, 19],
			[32, 8, 21], [33, 9, 20], [34, 10, 23], [35, 11, 22],
			[36, 44, 40], [37, 45, 41], [38, 46, 42], [39, 47, 43],
			[48, 52, 56], [49, 53, 57], [50, 54, 58], [51, 55, 59]]
	},
	Polyhedron{
		name:      'TruncatedDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.5
			z: 2.927051
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -2.927051
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 2.927051
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -2.927051
		}, Vertex{
			x: 2.927051
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 2.927051
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -2.927051
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -2.927051
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 2.927051
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -2.927051
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 2.927051
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -2.927051
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 2.618034
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: -2.618034
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 2.618034
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: -2.618034
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 2.618034
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: -2.618034
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 2.618034
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: -2.618034
		}, Vertex{
			x: 2.618034
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 2.618034
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 2.618034
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 2.618034
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: -2.618034
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: -2.618034
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: -2.618034
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: -2.618034
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 2.618034
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 2.618034
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: -2.618034
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: -2.618034
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 2.618034
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 2.618034
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: -2.618034
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: -2.618034
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: 1.618034
			z: 2.118034
		}, Vertex{
			x: 1.309017
			y: 1.618034
			z: -2.118034
		}, Vertex{
			x: 1.309017
			y: -1.618034
			z: 2.118034
		}, Vertex{
			x: 1.309017
			y: -1.618034
			z: -2.118034
		}, Vertex{
			x: -1.309017
			y: 1.618034
			z: 2.118034
		}, Vertex{
			x: -1.309017
			y: 1.618034
			z: -2.118034
		}, Vertex{
			x: -1.309017
			y: -1.618034
			z: 2.118034
		}, Vertex{
			x: -1.309017
			y: -1.618034
			z: -2.118034
		}, Vertex{
			x: 2.118034
			y: 1.309017
			z: 1.618034
		}, Vertex{
			x: 2.118034
			y: 1.309017
			z: -1.618034
		}, Vertex{
			x: 2.118034
			y: -1.309017
			z: 1.618034
		}, Vertex{
			x: 2.118034
			y: -1.309017
			z: -1.618034
		}, Vertex{
			x: -2.118034
			y: 1.309017
			z: 1.618034
		}, Vertex{
			x: -2.118034
			y: 1.309017
			z: -1.618034
		}, Vertex{
			x: -2.118034
			y: -1.309017
			z: 1.618034
		}, Vertex{
			x: -2.118034
			y: -1.309017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 2.118034
			z: 1.309017
		}, Vertex{
			x: 1.618034
			y: 2.118034
			z: -1.309017
		}, Vertex{
			x: 1.618034
			y: -2.118034
			z: 1.309017
		}, Vertex{
			x: 1.618034
			y: -2.118034
			z: -1.309017
		}, Vertex{
			x: -1.618034
			y: 2.118034
			z: 1.309017
		}, Vertex{
			x: -1.618034
			y: 2.118034
			z: -1.309017
		}, Vertex{
			x: -1.618034
			y: -2.118034
			z: 1.309017
		}, Vertex{
			x: -1.618034
			y: -2.118034
			z: -1.309017
		}]
		faces:     [[0, 2, 14, 38, 46, 22, 20, 44, 36, 12], [1, 3, 19, 43, 51, 27, 25, 49, 41, 17],
			[2, 0, 16, 40, 48, 24, 26, 50, 42, 18], [3, 1, 13, 37, 45, 21, 23, 47, 39, 15],
			[4, 5, 21, 45, 53, 29, 28, 52, 44, 20], [5, 4, 22, 46, 54, 30, 31, 55, 47, 23],
			[6, 7, 27, 51, 59, 35, 34, 58, 50, 26], [7, 6, 24, 48, 56, 32, 33, 57, 49, 25],
			[8, 10, 32, 56, 40, 16, 12, 36, 52, 28], [9, 11, 35, 59, 43, 19, 15, 39, 55, 31],
			[10, 8, 29, 53, 37, 13, 17, 41, 57, 33], [11, 9, 30, 54, 38, 14, 18, 42, 58, 34],
			[0, 12, 16], [1, 17, 13], [2, 18, 14], [3, 15, 19],
			[4, 20, 22], [5, 23, 21], [6, 26, 24], [7, 25, 27],
			[8, 28, 29], [9, 31, 30], [10, 33, 32], [11, 34, 35],
			[36, 44, 52], [37, 53, 45], [38, 54, 46], [39, 47, 55],
			[40, 56, 48], [41, 49, 57], [42, 50, 58], [43, 59, 51]]
	},
	Polyhedron{
		name:      'SmallDitrigonalDodecacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 2.427051
			y: 0.0
			z: 3.927051
		}, Vertex{
			x: 2.427051
			y: 0.0
			z: -3.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: 3.927051
		}, Vertex{
			x: -2.427051
			y: 0.0
			z: -3.927051
		}, Vertex{
			x: 3.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: 3.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: -3.927051
			y: 2.427051
			z: 0.0
		}, Vertex{
			x: -3.927051
			y: -2.427051
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 3.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: 3.927051
			z: -2.427051
		}, Vertex{
			x: 0.0
			y: -3.927051
			z: 2.427051
		}, Vertex{
			x: 0.0
			y: -3.927051
			z: -2.427051
		}, Vertex{
			x: 0.0
			y: 0.5970241
			z: 1.563030
		}, Vertex{
			x: 0.0
			y: 0.5970241
			z: -1.563030
		}, Vertex{
			x: 0.0
			y: -0.5970241
			z: 1.563030
		}, Vertex{
			x: 0.0
			y: -0.5970241
			z: -1.563030
		}, Vertex{
			x: 1.563030
			y: 0.0
			z: 0.5970241
		}, Vertex{
			x: 1.563030
			y: 0.0
			z: -0.5970241
		}, Vertex{
			x: -1.563030
			y: 0.0
			z: 0.5970241
		}, Vertex{
			x: -1.563030
			y: 0.0
			z: -0.5970241
		}, Vertex{
			x: 0.5970241
			y: 1.563030
			z: 0.0
		}, Vertex{
			x: 0.5970241
			y: -1.563030
			z: 0.0
		}, Vertex{
			x: -0.5970241
			y: 1.563030
			z: 0.0
		}, Vertex{
			x: -0.5970241
			y: -1.563030
			z: 0.0
		}, Vertex{
			x: 0.8702681
			y: 0.0
			z: 1.408123
		}, Vertex{
			x: 0.8702681
			y: 0.0
			z: -1.408123
		}, Vertex{
			x: -0.8702681
			y: 0.0
			z: 1.408123
		}, Vertex{
			x: -0.8702681
			y: 0.0
			z: -1.408123
		}, Vertex{
			x: 1.408123
			y: 0.8702681
			z: 0.0
		}, Vertex{
			x: 1.408123
			y: -0.8702681
			z: 0.0
		}, Vertex{
			x: -1.408123
			y: 0.8702681
			z: 0.0
		}, Vertex{
			x: -1.408123
			y: -0.8702681
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.408123
			z: 0.8702681
		}, Vertex{
			x: 0.0
			y: 1.408123
			z: -0.8702681
		}, Vertex{
			x: 0.0
			y: -1.408123
			z: 0.8702681
		}, Vertex{
			x: 0.0
			y: -1.408123
			z: -0.8702681
		}, Vertex{
			x: 0.9660054
			y: 0.9660054
			z: 0.9660054
		}, Vertex{
			x: 0.9660054
			y: 0.9660054
			z: -0.9660054
		}, Vertex{
			x: 0.9660054
			y: -0.9660054
			z: 0.9660054
		}, Vertex{
			x: 0.9660054
			y: -0.9660054
			z: -0.9660054
		}, Vertex{
			x: -0.9660054
			y: 0.9660054
			z: 0.9660054
		}, Vertex{
			x: -0.9660054
			y: 0.9660054
			z: -0.9660054
		}, Vertex{
			x: -0.9660054
			y: -0.9660054
			z: 0.9660054
		}, Vertex{
			x: -0.9660054
			y: -0.9660054
			z: -0.9660054
		}]
		faces:     [[24, 2, 38, 4], [24, 4, 12, 10], [24, 10, 16, 8],
			[24, 8, 14, 5], [24, 5, 36, 2], [25, 4, 39, 3], [25, 3, 37, 5],
			[25, 5, 15, 9], [25, 9, 17, 11], [25, 11, 13, 4],
			[26, 0, 40, 7], [26, 7, 14, 8], [26, 8, 18, 10], [26, 10, 12, 6],
			[26, 6, 42, 0], [27, 1, 43, 6], [27, 6, 13, 11], [27, 11, 19, 9],
			[27, 9, 15, 7], [27, 7, 41, 1], [28, 0, 17, 9], [28, 9, 36, 5],
			[28, 5, 37, 8], [28, 8, 16, 1], [28, 1, 20, 0], [29, 0, 21, 1],
			[29, 1, 16, 10], [29, 10, 39, 4], [29, 4, 38, 11],
			[29, 11, 17, 0], [30, 2, 22, 3], [30, 3, 18, 8], [30, 8, 41, 7],
			[30, 7, 40, 9], [30, 9, 19, 2], [31, 2, 19, 11], [31, 11, 42, 6],
			[31, 6, 43, 10], [31, 10, 18, 3], [31, 3, 23, 2],
			[32, 0, 20, 6], [32, 6, 12, 4], [32, 4, 22, 2], [32, 2, 36, 9],
			[32, 9, 40, 0], [33, 1, 41, 8], [33, 8, 37, 3], [33, 3, 22, 4],
			[33, 4, 13, 6], [33, 6, 20, 1], [34, 0, 42, 11], [34, 11, 38, 2],
			[34, 2, 23, 5], [34, 5, 14, 7], [34, 7, 21, 0], [35, 1, 21, 7],
			[35, 7, 15, 5], [35, 5, 23, 3], [35, 3, 39, 10], [35, 10, 43, 1]]
	},
	Polyhedron{
		name:      'InvertedSnubDodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.6760278
			y: 0.3626335
			z: 0.3698073
		}, Vertex{
			x: 0.6760278
			y: -0.3626335
			z: -0.3698073
		}, Vertex{
			x: -0.6760278
			y: -0.3626335
			z: 0.3698073
		}, Vertex{
			x: -0.6760278
			y: 0.3626335
			z: -0.3698073
		}, Vertex{
			x: 0.3698073
			y: 0.6760278
			z: 0.3626335
		}, Vertex{
			x: 0.3698073
			y: -0.6760278
			z: -0.3626335
		}, Vertex{
			x: -0.3698073
			y: -0.6760278
			z: 0.3626335
		}, Vertex{
			x: -0.3698073
			y: 0.6760278
			z: -0.3626335
		}, Vertex{
			x: 0.3626335
			y: 0.3698073
			z: 0.6760278
		}, Vertex{
			x: 0.3626335
			y: -0.3698073
			z: -0.6760278
		}, Vertex{
			x: -0.3626335
			y: -0.3698073
			z: 0.6760278
		}, Vertex{
			x: -0.3626335
			y: 0.3698073
			z: -0.6760278
		}, Vertex{
			x: 0.1589139
			y: 0.4740742
			z: 0.6894012
		}, Vertex{
			x: 0.1589139
			y: -0.4740742
			z: -0.6894012
		}, Vertex{
			x: -0.1589139
			y: -0.4740742
			z: 0.6894012
		}, Vertex{
			x: -0.1589139
			y: 0.4740742
			z: -0.6894012
		}, Vertex{
			x: 0.6894012
			y: -0.1589139
			z: -0.4740742
		}, Vertex{
			x: 0.6894012
			y: 0.1589139
			z: 0.4740742
		}, Vertex{
			x: -0.6894012
			y: 0.1589139
			z: -0.4740742
		}, Vertex{
			x: -0.6894012
			y: -0.1589139
			z: 0.4740742
		}, Vertex{
			x: -0.4740742
			y: -0.6894012
			z: 0.1589139
		}, Vertex{
			x: -0.4740742
			y: 0.6894012
			z: -0.1589139
		}, Vertex{
			x: 0.4740742
			y: 0.6894012
			z: 0.1589139
		}, Vertex{
			x: 0.4740742
			y: -0.6894012
			z: -0.1589139
		}, Vertex{
			x: -0.5171138
			y: 0.6197617
			z: 0.2715931
		}, Vertex{
			x: -0.5171138
			y: -0.6197617
			z: -0.2715931
		}, Vertex{
			x: 0.5171138
			y: -0.6197617
			z: 0.2715931
		}, Vertex{
			x: 0.5171138
			y: 0.6197617
			z: -0.2715931
		}, Vertex{
			x: 0.2715931
			y: -0.5171138
			z: 0.6197617
		}, Vertex{
			x: 0.2715931
			y: 0.5171138
			z: -0.6197617
		}, Vertex{
			x: -0.2715931
			y: 0.5171138
			z: 0.6197617
		}, Vertex{
			x: -0.2715931
			y: -0.5171138
			z: -0.6197617
		}, Vertex{
			x: 0.6197617
			y: 0.2715931
			z: -0.5171138
		}, Vertex{
			x: 0.6197617
			y: -0.2715931
			z: 0.5171138
		}, Vertex{
			x: -0.6197617
			y: -0.2715931
			z: -0.5171138
		}, Vertex{
			x: -0.6197617
			y: 0.2715931
			z: 0.5171138
		}, Vertex{
			x: 0.7456673
			y: -0.2499544
			z: 0.3267677
		}, Vertex{
			x: 0.7456673
			y: 0.2499544
			z: -0.3267677
		}, Vertex{
			x: -0.7456673
			y: 0.2499544
			z: 0.3267677
		}, Vertex{
			x: -0.7456673
			y: -0.2499544
			z: -0.3267677
		}, Vertex{
			x: 0.3267677
			y: 0.7456673
			z: -0.2499544
		}, Vertex{
			x: 0.3267677
			y: -0.7456673
			z: 0.2499544
		}, Vertex{
			x: -0.3267677
			y: -0.7456673
			z: -0.2499544
		}, Vertex{
			x: -0.3267677
			y: 0.7456673
			z: 0.2499544
		}, Vertex{
			x: -0.2499544
			y: 0.3267677
			z: 0.7456673
		}, Vertex{
			x: -0.2499544
			y: -0.3267677
			z: -0.7456673
		}, Vertex{
			x: 0.2499544
			y: -0.3267677
			z: 0.7456673
		}, Vertex{
			x: 0.2499544
			y: 0.3267677
			z: -0.7456673
		}, Vertex{
			x: -0.09104044
			y: -0.06963955
			z: 0.8438816
		}, Vertex{
			x: -0.09104044
			y: 0.06963955
			z: -0.8438816
		}, Vertex{
			x: 0.09104044
			y: 0.06963955
			z: 0.8438816
		}, Vertex{
			x: 0.09104044
			y: -0.06963955
			z: -0.8438816
		}, Vertex{
			x: 0.8438816
			y: 0.09104044
			z: 0.06963955
		}, Vertex{
			x: 0.8438816
			y: -0.09104044
			z: -0.06963955
		}, Vertex{
			x: -0.8438816
			y: -0.09104044
			z: 0.06963955
		}, Vertex{
			x: -0.8438816
			y: 0.09104044
			z: -0.06963955
		}, Vertex{
			x: 0.06963955
			y: -0.8438816
			z: -0.09104044
		}, Vertex{
			x: 0.06963955
			y: 0.8438816
			z: 0.09104044
		}, Vertex{
			x: -0.06963955
			y: 0.8438816
			z: -0.09104044
		}, Vertex{
			x: -0.06963955
			y: -0.8438816
			z: 0.09104044
		}]
		faces:     [[0, 28, 12, 36, 48], [1, 29, 13, 37, 49],
			[2, 30, 14, 38, 50], [3, 31, 15, 39, 51], [4, 32, 17, 40, 53],
			[5, 33, 16, 41, 52], [6, 34, 19, 42, 55], [7, 35, 18, 43, 54],
			[8, 24, 22, 44, 58], [9, 25, 23, 45, 59], [10, 26, 20, 46, 56],
			[11, 27, 21, 47, 57], [0, 26, 42, 18, 58], [1, 27, 43, 19, 59],
			[2, 24, 40, 16, 56], [3, 25, 41, 17, 57], [4, 29, 45, 20, 48],
			[5, 28, 44, 21, 49], [6, 31, 47, 22, 50], [7, 30, 46, 23, 51],
			[8, 35, 39, 13, 53], [9, 34, 38, 12, 52], [10, 33, 37, 15, 55],
			[11, 32, 36, 14, 54], [0, 58, 44], [1, 59, 45], [2, 56, 46],
			[3, 57, 47], [4, 48, 36], [5, 49, 37], [6, 50, 38],
			[7, 51, 39], [8, 53, 40], [9, 52, 41], [10, 55, 42],
			[11, 54, 43], [12, 38, 14], [13, 39, 15], [14, 36, 12],
			[15, 37, 13], [16, 40, 17], [17, 41, 16], [18, 42, 19],
			[19, 43, 18], [20, 45, 23], [21, 44, 22], [22, 47, 21],
			[23, 46, 20], [24, 2, 50], [25, 3, 51], [26, 0, 48],
			[27, 1, 49], [28, 5, 52], [29, 4, 53], [30, 7, 54],
			[31, 6, 55], [32, 11, 57], [33, 10, 56], [34, 9, 59],
			[35, 8, 58], [36, 32, 4], [37, 33, 5], [38, 34, 6],
			[39, 35, 7], [40, 24, 8], [41, 25, 9], [42, 26, 10],
			[43, 27, 11], [44, 28, 0], [45, 29, 1], [46, 30, 2],
			[47, 31, 3], [48, 20, 26], [49, 21, 27], [50, 22, 24],
			[51, 23, 25], [52, 12, 28], [53, 13, 29], [54, 14, 30],
			[55, 15, 31], [56, 16, 33], [57, 17, 32], [58, 18, 35],
			[59, 19, 34]]
	},
	Polyhedron{
		name:      'StellatedTruncatedHexahedron'
		vertexes_: [Vertex{
			x: -0.2071068
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: -0.2071068
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: 0.2071068
		}]
		faces:     [[0, 2, 10, 11, 3, 1, 9, 8], [0, 16, 20, 4, 6, 22, 18, 2],
			[12, 13, 5, 7, 15, 14, 6, 4], [12, 20, 16, 8, 9, 17, 21, 13],
			[19, 23, 7, 5, 21, 17, 1, 3], [19, 11, 10, 18, 22, 14, 15, 23],
			[0, 8, 16], [1, 17, 9], [2, 18, 10], [3, 11, 19],
			[4, 20, 12], [5, 13, 21], [6, 14, 22], [7, 23, 15]]
	},
	Polyhedron{
		name:      'GreatTriakisOctahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: -0.4142136
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 0.4142136
		}, Vertex{
			x: -0.4142136
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.4142136
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.4142136
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.4142136
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[6, 0, 2], [6, 2, 4], [6, 4, 0], [7, 1, 4],
			[7, 4, 2], [7, 2, 1], [8, 0, 5], [8, 5, 2], [8, 2, 0],
			[9, 1, 2], [9, 2, 5], [9, 5, 1], [10, 0, 4], [10, 4, 3],
			[10, 3, 0], [11, 1, 3], [11, 3, 4], [11, 4, 1], [12, 0, 3],
			[12, 3, 5], [12, 5, 0], [13, 1, 5], [13, 5, 3], [13, 3, 1]]
	},
	Polyhedron{
		name:      'DeltoidalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 2.236068
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -2.236068
		}, Vertex{
			x: 2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -2.236068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.236068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -2.236068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7834576
			z: 2.051119
		}, Vertex{
			x: 0.0
			y: 0.7834576
			z: -2.051119
		}, Vertex{
			x: 0.0
			y: -0.7834576
			z: 2.051119
		}, Vertex{
			x: 0.0
			y: -0.7834576
			z: -2.051119
		}, Vertex{
			x: 2.051119
			y: 0.0
			z: 0.7834576
		}, Vertex{
			x: 2.051119
			y: 0.0
			z: -0.7834576
		}, Vertex{
			x: -2.051119
			y: 0.0
			z: 0.7834576
		}, Vertex{
			x: -2.051119
			y: 0.0
			z: -0.7834576
		}, Vertex{
			x: 0.7834576
			y: 2.051119
			z: 0.0
		}, Vertex{
			x: 0.7834576
			y: -2.051119
			z: 0.0
		}, Vertex{
			x: -0.7834576
			y: 2.051119
			z: 0.0
		}, Vertex{
			x: -0.7834576
			y: -2.051119
			z: 0.0
		}, Vertex{
			x: 1.206011
			y: 0.0
			z: 1.951367
		}, Vertex{
			x: 1.206011
			y: 0.0
			z: -1.951367
		}, Vertex{
			x: -1.206011
			y: 0.0
			z: 1.951367
		}, Vertex{
			x: -1.206011
			y: 0.0
			z: -1.951367
		}, Vertex{
			x: 1.951367
			y: 1.206011
			z: 0.0
		}, Vertex{
			x: 1.951367
			y: -1.206011
			z: 0.0
		}, Vertex{
			x: -1.951367
			y: 1.206011
			z: 0.0
		}, Vertex{
			x: -1.951367
			y: -1.206011
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.951367
			z: 1.206011
		}, Vertex{
			x: 0.0
			y: 1.951367
			z: -1.206011
		}, Vertex{
			x: 0.0
			y: -1.951367
			z: 1.206011
		}, Vertex{
			x: 0.0
			y: -1.951367
			z: -1.206011
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: 0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: 1.118034
			z: -1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: 1.809017
		}, Vertex{
			x: -0.690983
			y: -1.118034
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: 1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: 1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: 0.690983
			z: -1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: 1.118034
		}, Vertex{
			x: -1.809017
			y: -0.690983
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: 1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: 1.809017
			z: -0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: 0.690983
		}, Vertex{
			x: -1.118034
			y: -1.809017
			z: -0.690983
		}, Vertex{
			x: 1.267661
			y: 1.267661
			z: 1.267661
		}, Vertex{
			x: 1.267661
			y: 1.267661
			z: -1.267661
		}, Vertex{
			x: 1.267661
			y: -1.267661
			z: 1.267661
		}, Vertex{
			x: 1.267661
			y: -1.267661
			z: -1.267661
		}, Vertex{
			x: -1.267661
			y: 1.267661
			z: 1.267661
		}, Vertex{
			x: -1.267661
			y: 1.267661
			z: -1.267661
		}, Vertex{
			x: -1.267661
			y: -1.267661
			z: 1.267661
		}, Vertex{
			x: -1.267661
			y: -1.267661
			z: -1.267661
		}]
		faces:     [[18, 0, 8, 32], [18, 32, 56, 40], [18, 40, 10, 38],
			[18, 38, 54, 30], [18, 30, 6, 0], [19, 1, 7, 31],
			[19, 31, 55, 39], [19, 39, 11, 41], [19, 41, 57, 33],
			[19, 33, 9, 1], [20, 0, 6, 34], [20, 34, 58, 42],
			[20, 42, 12, 44], [20, 44, 60, 36], [20, 36, 8, 0],
			[21, 1, 9, 37], [21, 37, 61, 45], [21, 45, 13, 43],
			[21, 43, 59, 35], [21, 35, 7, 1], [22, 2, 11, 39],
			[22, 39, 55, 47], [22, 47, 14, 46], [22, 46, 54, 38],
			[22, 38, 10, 2], [23, 2, 10, 40], [23, 40, 56, 48],
			[23, 48, 15, 49], [23, 49, 57, 41], [23, 41, 11, 2],
			[24, 3, 12, 42], [24, 42, 58, 50], [24, 50, 16, 51],
			[24, 51, 59, 43], [24, 43, 13, 3], [25, 3, 13, 45],
			[25, 45, 61, 53], [25, 53, 17, 52], [25, 52, 60, 44],
			[25, 44, 12, 3], [26, 4, 16, 50], [26, 50, 58, 34],
			[26, 34, 6, 30], [26, 30, 54, 46], [26, 46, 14, 4],
			[27, 4, 14, 47], [27, 47, 55, 31], [27, 31, 7, 35],
			[27, 35, 59, 51], [27, 51, 16, 4], [28, 5, 15, 48],
			[28, 48, 56, 32], [28, 32, 8, 36], [28, 36, 60, 52],
			[28, 52, 17, 5], [29, 5, 17, 53], [29, 53, 61, 37],
			[29, 37, 9, 33], [29, 33, 57, 49], [29, 49, 15, 5]]
	},
	Polyhedron{
		name:      'MedialInvertedPentagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.6034342
			z: -0.3729428
		}, Vertex{
			x: 0.0
			y: 0.6034342
			z: 0.3729428
		}, Vertex{
			x: 0.0
			y: -0.6034342
			z: -0.3729428
		}, Vertex{
			x: 0.0
			y: -0.6034342
			z: 0.3729428
		}, Vertex{
			x: 0.6034342
			y: -0.3729428
			z: 0.0
		}, Vertex{
			x: -0.6034342
			y: -0.3729428
			z: 0.0
		}, Vertex{
			x: 0.6034342
			y: 0.3729428
			z: 0.0
		}, Vertex{
			x: -0.6034342
			y: 0.3729428
			z: 0.0
		}, Vertex{
			x: -0.3729428
			y: 0.0
			z: 0.6034342
		}, Vertex{
			x: -0.3729428
			y: 0.0
			z: -0.6034342
		}, Vertex{
			x: 0.3729428
			y: 0.0
			z: 0.6034342
		}, Vertex{
			x: 0.3729428
			y: 0.0
			z: -0.6034342
		}, Vertex{
			x: 0.301403
			y: 0.1010330
			z: 0.6894012
		}, Vertex{
			x: -0.301403
			y: 0.1010330
			z: -0.6894012
		}, Vertex{
			x: -0.301403
			y: -0.1010330
			z: 0.6894012
		}, Vertex{
			x: 0.301403
			y: -0.1010330
			z: -0.6894012
		}, Vertex{
			x: -0.1010330
			y: 0.6894012
			z: -0.301403
		}, Vertex{
			x: 0.1010330
			y: 0.6894012
			z: 0.301403
		}, Vertex{
			x: 0.1010330
			y: -0.6894012
			z: -0.301403
		}, Vertex{
			x: -0.1010330
			y: -0.6894012
			z: 0.301403
		}, Vertex{
			x: -0.6894012
			y: -0.301403
			z: 0.1010330
		}, Vertex{
			x: 0.6894012
			y: -0.301403
			z: -0.1010330
		}, Vertex{
			x: 0.6894012
			y: 0.301403
			z: 0.1010330
		}, Vertex{
			x: -0.6894012
			y: 0.301403
			z: -0.1010330
		}, Vertex{
			x: 0.1320814
			y: -0.6003594
			z: -0.4454756
		}, Vertex{
			x: -0.1320814
			y: -0.6003594
			z: 0.4454756
		}, Vertex{
			x: -0.1320814
			y: 0.6003594
			z: -0.4454756
		}, Vertex{
			x: 0.1320814
			y: 0.6003594
			z: 0.4454756
		}, Vertex{
			x: -0.6003594
			y: -0.4454756
			z: 0.1320814
		}, Vertex{
			x: 0.6003594
			y: -0.4454756
			z: -0.1320814
		}, Vertex{
			x: 0.6003594
			y: 0.4454756
			z: 0.1320814
		}, Vertex{
			x: -0.6003594
			y: 0.4454756
			z: -0.1320814
		}, Vertex{
			x: -0.4454756
			y: 0.1320814
			z: -0.6003594
		}, Vertex{
			x: 0.4454756
			y: 0.1320814
			z: 0.6003594
		}, Vertex{
			x: 0.4454756
			y: -0.1320814
			z: -0.6003594
		}, Vertex{
			x: -0.4454756
			y: -0.1320814
			z: 0.6003594
		}, Vertex{
			x: 0.0
			y: 9.901372
			z: -6.119384
		}, Vertex{
			x: 0.0
			y: 9.901372
			z: 6.119384
		}, Vertex{
			x: 0.0
			y: -9.901372
			z: -6.119384
		}, Vertex{
			x: 0.0
			y: -9.901372
			z: 6.119384
		}, Vertex{
			x: 9.901372
			y: -6.119384
			z: 0.0
		}, Vertex{
			x: -9.901372
			y: -6.119384
			z: 0.0
		}, Vertex{
			x: 9.901372
			y: 6.119384
			z: 0.0
		}, Vertex{
			x: -9.901372
			y: 6.119384
			z: 0.0
		}, Vertex{
			x: -6.119384
			y: 0.0
			z: 9.901372
		}, Vertex{
			x: -6.119384
			y: 0.0
			z: -9.901372
		}, Vertex{
			x: 6.119384
			y: 0.0
			z: 9.901372
		}, Vertex{
			x: 6.119384
			y: 0.0
			z: -9.901372
		}, Vertex{
			x: -0.06963955
			y: -0.7013925
			z: -0.2820008
		}, Vertex{
			x: 0.06963955
			y: -0.7013925
			z: 0.2820008
		}, Vertex{
			x: 0.06963955
			y: 0.7013925
			z: -0.2820008
		}, Vertex{
			x: -0.06963955
			y: 0.7013925
			z: 0.2820008
		}, Vertex{
			x: 0.7013925
			y: -0.2820008
			z: 0.06963955
		}, Vertex{
			x: -0.7013925
			y: -0.2820008
			z: -0.06963955
		}, Vertex{
			x: -0.7013925
			y: 0.2820008
			z: 0.06963955
		}, Vertex{
			x: 0.7013925
			y: 0.2820008
			z: -0.06963955
		}, Vertex{
			x: 0.2820008
			y: 0.06963955
			z: -0.7013925
		}, Vertex{
			x: -0.2820008
			y: 0.06963955
			z: 0.7013925
		}, Vertex{
			x: -0.2820008
			y: -0.06963955
			z: -0.7013925
		}, Vertex{
			x: 0.2820008
			y: -0.06963955
			z: 0.7013925
		}, Vertex{
			x: -0.6197617
			y: -0.4140822
			z: -0.1440726
		}, Vertex{
			x: 0.6197617
			y: -0.4140822
			z: 0.1440726
		}, Vertex{
			x: 0.6197617
			y: 0.4140822
			z: -0.1440726
		}, Vertex{
			x: -0.6197617
			y: 0.4140822
			z: 0.1440726
		}, Vertex{
			x: 0.4140822
			y: -0.1440726
			z: 0.6197617
		}, Vertex{
			x: -0.4140822
			y: -0.1440726
			z: -0.6197617
		}, Vertex{
			x: -0.4140822
			y: 0.1440726
			z: 0.6197617
		}, Vertex{
			x: 0.4140822
			y: 0.1440726
			z: -0.6197617
		}, Vertex{
			x: 0.1440726
			y: 0.6197617
			z: -0.4140822
		}, Vertex{
			x: -0.1440726
			y: 0.6197617
			z: 0.4140822
		}, Vertex{
			x: -0.1440726
			y: -0.6197617
			z: -0.4140822
		}, Vertex{
			x: 0.1440726
			y: -0.6197617
			z: 0.4140822
		}, Vertex{
			x: -0.5151151
			y: 0.01940221
			z: 0.5573198
		}, Vertex{
			x: 0.5151151
			y: 0.01940221
			z: -0.5573198
		}, Vertex{
			x: 0.5151151
			y: -0.01940221
			z: 0.5573198
		}, Vertex{
			x: -0.5151151
			y: -0.01940221
			z: -0.5573198
		}, Vertex{
			x: 0.01940221
			y: 0.5573198
			z: -0.5151151
		}, Vertex{
			x: -0.01940221
			y: 0.5573198
			z: 0.5151151
		}, Vertex{
			x: -0.01940221
			y: -0.5573198
			z: -0.5151151
		}, Vertex{
			x: 0.01940221
			y: -0.5573198
			z: 0.5151151
		}, Vertex{
			x: 0.5573198
			y: -0.5151151
			z: 0.01940221
		}, Vertex{
			x: -0.5573198
			y: -0.5151151
			z: -0.01940221
		}, Vertex{
			x: -0.5573198
			y: 0.5151151
			z: 0.01940221
		}, Vertex{
			x: 0.5573198
			y: 0.5151151
			z: -0.01940221
		}]
		faces:     [[0, 16, 17, 40, 76], [0, 76, 32, 44, 50],
			[0, 50, 62, 38, 26], [0, 26, 82, 46, 68], [0, 68, 56, 41, 16],
			[1, 17, 16, 41, 77], [1, 77, 33, 47, 51], [1, 51, 63, 39, 27],
			[1, 27, 83, 45, 69], [1, 69, 57, 40, 17], [2, 18, 19, 43, 78],
			[2, 78, 34, 46, 48], [2, 48, 60, 36, 24], [2, 24, 80, 44, 70],
			[2, 70, 58, 42, 18], [3, 19, 18, 42, 79], [3, 79, 35, 45, 49],
			[3, 49, 61, 37, 25], [3, 25, 81, 47, 71], [3, 71, 59, 43, 19],
			[4, 21, 22, 44, 80], [4, 80, 24, 36, 52], [4, 52, 64, 41, 29],
			[4, 29, 73, 37, 61], [4, 61, 49, 45, 21], [5, 20, 23, 47, 81],
			[5, 81, 25, 37, 53], [5, 53, 65, 40, 28], [5, 28, 72, 36, 60],
			[5, 60, 48, 46, 20], [6, 22, 21, 45, 83], [6, 83, 27, 39, 55],
			[6, 55, 67, 43, 30], [6, 30, 74, 38, 62], [6, 62, 50, 44, 22],
			[7, 23, 20, 46, 82], [7, 82, 26, 38, 54], [7, 54, 66, 42, 31],
			[7, 31, 75, 39, 63], [7, 63, 51, 47, 23], [8, 14, 12, 36, 72],
			[8, 72, 28, 40, 57], [8, 57, 69, 45, 35], [8, 35, 79, 42, 66],
			[8, 66, 54, 38, 14], [9, 13, 15, 39, 75], [9, 75, 31, 42, 58],
			[9, 58, 70, 44, 32], [9, 32, 76, 40, 65], [9, 65, 53, 37, 13],
			[10, 12, 14, 38, 74], [10, 74, 30, 43, 59], [10, 59, 71, 47, 33],
			[10, 33, 77, 41, 64], [10, 64, 52, 36, 12], [11, 15, 13, 37, 73],
			[11, 73, 29, 41, 56], [11, 56, 68, 46, 34], [11, 34, 78, 43, 67],
			[11, 67, 55, 39, 15]]
	},
	Polyhedron{
		name:      'SmallDodecicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: 2.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 2.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: -0.5
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: 1.618034
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: -1.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: 1.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: -1.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: 1.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: -1.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: 1.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: 1.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: 1.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: 1.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: -1.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: -1.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: -1.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: -1.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: 1.618034
			z: -1.309017
		}, Vertex{
			x: 0.809017
			y: -1.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: -1.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: 1.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: 1.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: -1.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: -1.618034
			z: -1.309017
		}]
		faces:     [[0, 24, 56, 48, 12, 14, 50, 58, 26, 2], [0, 36, 44, 32, 17, 21, 34, 48, 40,
			4],
			[7, 3, 39, 47, 33, 18, 22, 35, 51, 43], [7, 5, 25, 53, 45, 9, 11, 47, 55, 27],
			[10, 8, 44, 52, 24, 4, 6, 26, 54, 46], [10, 11, 29, 37, 53, 17, 16, 52, 36, 28],
			[13, 31, 43, 59, 23, 22, 58, 42, 30, 12], [13, 49, 57, 25, 1, 3, 27, 59, 51, 15],
			[19, 33, 46, 38, 2, 6, 42, 50, 35, 23], [19, 55, 39, 29, 9, 8, 28, 38, 54, 18],
			[20, 16, 32, 45, 37, 1, 5, 41, 49, 34], [20, 21, 57, 41, 31, 15, 14, 30, 40, 56],
			[24, 52, 16, 20, 56], [25, 57, 21, 17, 53], [26, 58, 22, 18, 54],
			[27, 55, 19, 23, 59], [28, 36, 0, 2, 38], [29, 39, 3, 1, 37],
			[30, 42, 6, 4, 40], [31, 41, 5, 7, 43], [32, 44, 8, 9, 45],
			[33, 47, 11, 10, 46], [34, 49, 13, 12, 48], [35, 50, 14, 15, 51],
			[24, 0, 4], [25, 5, 1], [26, 6, 2], [27, 3, 7], [28, 8, 10],
			[29, 11, 9], [30, 14, 12], [31, 13, 15], [32, 16, 17],
			[33, 19, 18], [34, 21, 20], [35, 22, 23], [36, 52, 44],
			[37, 45, 53], [38, 46, 54], [39, 55, 47], [40, 48, 56],
			[41, 57, 49], [42, 58, 50], [43, 51, 59]]
	},
	Polyhedron{
		name:      'RhombicTriacontahedron'
		vertexes_: [Vertex{
			x: 0.9045085
			y: 0.0
			z: 1.463526
		}, Vertex{
			x: 0.9045085
			y: 0.0
			z: -1.463526
		}, Vertex{
			x: -0.9045085
			y: 0.0
			z: 1.463526
		}, Vertex{
			x: -0.9045085
			y: 0.0
			z: -1.463526
		}, Vertex{
			x: 1.463526
			y: 0.9045085
			z: 0.0
		}, Vertex{
			x: 1.463526
			y: -0.9045085
			z: 0.0
		}, Vertex{
			x: -1.463526
			y: 0.9045085
			z: 0.0
		}, Vertex{
			x: -1.463526
			y: -0.9045085
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.463526
			z: 0.9045085
		}, Vertex{
			x: 0.0
			y: 1.463526
			z: -0.9045085
		}, Vertex{
			x: 0.0
			y: -1.463526
			z: 0.9045085
		}, Vertex{
			x: 0.0
			y: -1.463526
			z: -0.9045085
		}, Vertex{
			x: 0.0
			y: 0.559017
			z: 1.463526
		}, Vertex{
			x: 0.0
			y: 0.559017
			z: -1.463526
		}, Vertex{
			x: 0.0
			y: -0.559017
			z: 1.463526
		}, Vertex{
			x: 0.0
			y: -0.559017
			z: -1.463526
		}, Vertex{
			x: 1.463526
			y: 0.0
			z: 0.559017
		}, Vertex{
			x: 1.463526
			y: 0.0
			z: -0.559017
		}, Vertex{
			x: -1.463526
			y: 0.0
			z: 0.559017
		}, Vertex{
			x: -1.463526
			y: 0.0
			z: -0.559017
		}, Vertex{
			x: 0.559017
			y: 1.463526
			z: 0.0
		}, Vertex{
			x: 0.559017
			y: -1.463526
			z: 0.0
		}, Vertex{
			x: -0.559017
			y: 1.463526
			z: 0.0
		}, Vertex{
			x: -0.559017
			y: -1.463526
			z: 0.0
		}, Vertex{
			x: 0.9045085
			y: 0.9045085
			z: 0.9045085
		}, Vertex{
			x: 0.9045085
			y: 0.9045085
			z: -0.9045085
		}, Vertex{
			x: 0.9045085
			y: -0.9045085
			z: 0.9045085
		}, Vertex{
			x: 0.9045085
			y: -0.9045085
			z: -0.9045085
		}, Vertex{
			x: -0.9045085
			y: 0.9045085
			z: 0.9045085
		}, Vertex{
			x: -0.9045085
			y: 0.9045085
			z: -0.9045085
		}, Vertex{
			x: -0.9045085
			y: -0.9045085
			z: 0.9045085
		}, Vertex{
			x: -0.9045085
			y: -0.9045085
			z: -0.9045085
		}]
		faces:     [[0, 12, 2, 14], [0, 14, 10, 26], [0, 26, 5, 16],
			[1, 13, 9, 25], [1, 25, 4, 17], [1, 17, 5, 27], [2, 28, 6, 18],
			[2, 18, 7, 30], [2, 30, 10, 14], [3, 19, 6, 29], [3, 29, 9, 13],
			[3, 13, 1, 15], [4, 20, 8, 24], [4, 24, 0, 16], [4, 16, 5, 17],
			[7, 18, 6, 19], [7, 19, 3, 31], [7, 31, 11, 23], [8, 22, 6, 28],
			[8, 28, 2, 12], [8, 12, 0, 24], [9, 29, 6, 22], [9, 22, 8, 20],
			[9, 20, 4, 25], [10, 30, 7, 23], [10, 23, 11, 21],
			[10, 21, 5, 26], [11, 31, 3, 15], [11, 15, 1, 27],
			[11, 27, 5, 21]]
	},
	Polyhedron{
		name:      'Dodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: -0.809017
		}]
		faces:     [[0, 2, 14, 4, 12], [0, 12, 8, 10, 16], [0, 16, 6, 18, 2],
			[7, 6, 16, 10, 17], [7, 17, 1, 3, 19], [7, 19, 11, 18, 6],
			[9, 11, 19, 3, 15], [9, 15, 5, 4, 14], [9, 14, 2, 18, 11],
			[13, 1, 17, 10, 8], [13, 8, 12, 4, 5], [13, 5, 15, 3, 1]]
	},
	Polyhedron{
		name:      'SmallIcosacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -1.809017
		}, Vertex{
			x: 0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.408123
			z: 0.8702681
		}, Vertex{
			x: 0.0
			y: -1.408123
			z: -0.8702681
		}, Vertex{
			x: 0.0
			y: 1.408123
			z: 0.8702681
		}, Vertex{
			x: 0.0
			y: 1.408123
			z: -0.8702681
		}, Vertex{
			x: -1.408123
			y: 0.8702681
			z: 0.0
		}, Vertex{
			x: 1.408123
			y: 0.8702681
			z: 0.0
		}, Vertex{
			x: -1.408123
			y: -0.8702681
			z: 0.0
		}, Vertex{
			x: 1.408123
			y: -0.8702681
			z: 0.0
		}, Vertex{
			x: 0.8702681
			y: 0.0
			z: -1.408123
		}, Vertex{
			x: 0.8702681
			y: 0.0
			z: 1.408123
		}, Vertex{
			x: -0.8702681
			y: 0.0
			z: -1.408123
		}, Vertex{
			x: -0.8702681
			y: 0.0
			z: 1.408123
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: -1.563030
			y: 0.0
			z: -0.5970241
		}, Vertex{
			x: -1.563030
			y: 0.0
			z: 0.5970241
		}, Vertex{
			x: 1.563030
			y: 0.0
			z: -0.5970241
		}, Vertex{
			x: 1.563030
			y: 0.0
			z: 0.5970241
		}, Vertex{
			x: 0.0
			y: -0.5970241
			z: -1.563030
		}, Vertex{
			x: 0.0
			y: -0.5970241
			z: 1.563030
		}, Vertex{
			x: 0.0
			y: 0.5970241
			z: -1.563030
		}, Vertex{
			x: 0.0
			y: 0.5970241
			z: 1.563030
		}, Vertex{
			x: -0.5970241
			y: -1.563030
			z: 0.0
		}, Vertex{
			x: 0.5970241
			y: -1.563030
			z: 0.0
		}, Vertex{
			x: -0.5970241
			y: 1.563030
			z: 0.0
		}, Vertex{
			x: 0.5970241
			y: 1.563030
			z: 0.0
		}, Vertex{
			x: 0.9660054
			y: 0.9660054
			z: 0.9660054
		}, Vertex{
			x: 0.9660054
			y: 0.9660054
			z: -0.9660054
		}, Vertex{
			x: -0.9660054
			y: 0.9660054
			z: 0.9660054
		}, Vertex{
			x: -0.9660054
			y: 0.9660054
			z: -0.9660054
		}, Vertex{
			x: 0.9660054
			y: -0.9660054
			z: 0.9660054
		}, Vertex{
			x: 0.9660054
			y: -0.9660054
			z: -0.9660054
		}, Vertex{
			x: -0.9660054
			y: -0.9660054
			z: 0.9660054
		}, Vertex{
			x: -0.9660054
			y: -0.9660054
			z: -0.9660054
		}]
		faces:     [[12, 6, 50, 11], [12, 11, 41, 27], [12, 27, 37, 25],
			[12, 25, 40, 10], [12, 10, 48, 6], [13, 7, 49, 10],
			[13, 10, 40, 24], [13, 24, 36, 26], [13, 26, 41, 11],
			[13, 11, 51, 7], [14, 4, 44, 8], [14, 8, 42, 29],
			[14, 29, 39, 31], [14, 31, 43, 9], [14, 9, 46, 4],
			[15, 5, 47, 9], [15, 9, 43, 30], [15, 30, 38, 28],
			[15, 28, 42, 8], [15, 8, 45, 5], [16, 2, 46, 9], [16, 9, 47, 3],
			[16, 3, 33, 29], [16, 29, 42, 28], [16, 28, 32, 2],
			[17, 0, 34, 30], [17, 30, 43, 31], [17, 31, 35, 1],
			[17, 1, 45, 8], [17, 8, 44, 0], [18, 2, 32, 24], [18, 24, 40, 25],
			[18, 25, 33, 3], [18, 3, 51, 11], [18, 11, 50, 2],
			[19, 0, 48, 10], [19, 10, 49, 1], [19, 1, 35, 27],
			[19, 27, 41, 26], [19, 26, 34, 0], [20, 1, 49, 7],
			[20, 7, 38, 30], [20, 30, 34, 26], [20, 26, 36, 5],
			[20, 5, 45, 1], [21, 0, 44, 4], [21, 4, 37, 27], [21, 27, 35, 31],
			[21, 31, 39, 6], [21, 6, 48, 0], [22, 3, 47, 5], [22, 5, 36, 24],
			[22, 24, 32, 28], [22, 28, 38, 7], [22, 7, 51, 3],
			[23, 2, 50, 6], [23, 6, 39, 29], [23, 29, 33, 25],
			[23, 25, 37, 4], [23, 4, 46, 2]]
	},
	Polyhedron{
		name:      'Tetrahemihexahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: 0.0
		}]
		faces:     [[0, 2, 1, 3], [0, 5, 1, 4], [2, 4, 3, 5],
			[0, 2, 4], [0, 3, 5], [1, 2, 5], [1, 3, 4]]
	},
	Polyhedron{
		name:      'GreatIcosidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: -0.309017
			z: 0.5
		}]
		faces:     [[0, 8, 16, 14, 6], [0, 10, 18, 20, 12], [1, 7, 15, 17, 9],
			[1, 13, 21, 19, 11], [2, 15, 23, 22, 14], [2, 16, 24, 25, 17],
			[3, 18, 26, 27, 19], [3, 21, 29, 28, 20], [4, 23, 7, 11, 27],
			[4, 26, 10, 6, 22], [5, 24, 8, 12, 28], [5, 29, 13, 9, 25],
			[0, 6, 10], [0, 12, 8], [1, 9, 13], [1, 11, 7], [2, 14, 16],
			[2, 17, 15], [3, 19, 21], [3, 20, 18], [4, 22, 23],
			[4, 27, 26], [5, 25, 24], [5, 28, 29], [6, 14, 22],
			[7, 23, 15], [8, 24, 16], [9, 17, 25], [10, 26, 18],
			[11, 19, 27], [12, 20, 28], [13, 29, 21]]
	},
	Polyhedron{
		name:      'GreatSnubIcosidodecahedron'
		vertexes_: [Vertex{
			x: -0.3710472
			y: 0.3351477
			z: -0.6449711
		}, Vertex{
			x: 0.3710472
			y: 0.3351477
			z: 0.6449711
		}, Vertex{
			x: 0.3710472
			y: -0.3351477
			z: -0.6449711
		}, Vertex{
			x: -0.3710472
			y: -0.3351477
			z: 0.6449711
		}, Vertex{
			x: 0.3351477
			y: -0.6449711
			z: -0.3710472
		}, Vertex{
			x: -0.3351477
			y: -0.6449711
			z: 0.3710472
		}, Vertex{
			x: -0.3351477
			y: 0.6449711
			z: -0.3710472
		}, Vertex{
			x: 0.3351477
			y: 0.6449711
			z: 0.3710472
		}, Vertex{
			x: -0.6449711
			y: -0.3710472
			z: 0.3351477
		}, Vertex{
			x: 0.6449711
			y: -0.3710472
			z: -0.3351477
		}, Vertex{
			x: 0.6449711
			y: 0.3710472
			z: 0.3351477
		}, Vertex{
			x: -0.6449711
			y: 0.3710472
			z: -0.3351477
		}, Vertex{
			x: 0.5191027
			y: 0.5747065
			z: -0.2573568
		}, Vertex{
			x: -0.5191027
			y: 0.5747065
			z: 0.2573568
		}, Vertex{
			x: -0.5191027
			y: -0.5747065
			z: -0.2573568
		}, Vertex{
			x: 0.5191027
			y: -0.5747065
			z: 0.2573568
		}, Vertex{
			x: -0.5747065
			y: -0.2573568
			z: -0.5191027
		}, Vertex{
			x: 0.5747065
			y: -0.2573568
			z: 0.5191027
		}, Vertex{
			x: 0.5747065
			y: 0.2573568
			z: -0.5191027
		}, Vertex{
			x: -0.5747065
			y: 0.2573568
			z: 0.5191027
		}, Vertex{
			x: 0.2573568
			y: -0.5191027
			z: 0.5747065
		}, Vertex{
			x: -0.2573568
			y: -0.5191027
			z: -0.5747065
		}, Vertex{
			x: -0.2573568
			y: 0.5191027
			z: 0.5747065
		}, Vertex{
			x: 0.2573568
			y: 0.5191027
			z: -0.5747065
		}, Vertex{
			x: -0.7262353
			y: 0.2395588
			z: 0.2849236
		}, Vertex{
			x: 0.7262353
			y: 0.2395588
			z: -0.2849236
		}, Vertex{
			x: 0.7262353
			y: -0.2395588
			z: 0.2849236
		}, Vertex{
			x: -0.7262353
			y: -0.2395588
			z: -0.2849236
		}, Vertex{
			x: 0.2395588
			y: 0.2849236
			z: -0.7262353
		}, Vertex{
			x: -0.2395588
			y: 0.2849236
			z: 0.7262353
		}, Vertex{
			x: -0.2395588
			y: -0.2849236
			z: -0.7262353
		}, Vertex{
			x: 0.2395588
			y: -0.2849236
			z: 0.7262353
		}, Vertex{
			x: 0.2849236
			y: -0.7262353
			z: 0.2395588
		}, Vertex{
			x: -0.2849236
			y: -0.7262353
			z: -0.2395588
		}, Vertex{
			x: -0.2849236
			y: 0.7262353
			z: 0.2395588
		}, Vertex{
			x: 0.2849236
			y: 0.7262353
			z: -0.2395588
		}, Vertex{
			x: 0.08126428
			y: 0.8040263
			z: 0.1136904
		}, Vertex{
			x: -0.08126428
			y: 0.8040263
			z: -0.1136904
		}, Vertex{
			x: -0.08126428
			y: -0.8040263
			z: 0.1136904
		}, Vertex{
			x: 0.08126428
			y: -0.8040263
			z: -0.1136904
		}, Vertex{
			x: 0.8040263
			y: 0.1136904
			z: 0.08126428
		}, Vertex{
			x: -0.8040263
			y: 0.1136904
			z: -0.08126428
		}, Vertex{
			x: -0.8040263
			y: -0.1136904
			z: 0.08126428
		}, Vertex{
			x: 0.8040263
			y: -0.1136904
			z: -0.08126428
		}, Vertex{
			x: 0.1136904
			y: 0.08126428
			z: 0.8040263
		}, Vertex{
			x: -0.1136904
			y: 0.08126428
			z: -0.8040263
		}, Vertex{
			x: -0.1136904
			y: -0.08126428
			z: 0.8040263
		}, Vertex{
			x: 0.1136904
			y: -0.08126428
			z: -0.8040263
		}, Vertex{
			x: -0.4688786
			y: 0.6559708
			z: -0.1258684
		}, Vertex{
			x: 0.4688786
			y: 0.6559708
			z: 0.1258684
		}, Vertex{
			x: 0.4688786
			y: -0.6559708
			z: -0.1258684
		}, Vertex{
			x: -0.4688786
			y: -0.6559708
			z: 0.1258684
		}, Vertex{
			x: -0.6559708
			y: -0.1258684
			z: 0.4688786
		}, Vertex{
			x: 0.6559708
			y: -0.1258684
			z: -0.4688786
		}, Vertex{
			x: 0.6559708
			y: 0.1258684
			z: 0.4688786
		}, Vertex{
			x: -0.6559708
			y: 0.1258684
			z: -0.4688786
		}, Vertex{
			x: 0.1258684
			y: 0.4688786
			z: 0.6559708
		}, Vertex{
			x: -0.1258684
			y: 0.4688786
			z: -0.6559708
		}, Vertex{
			x: -0.1258684
			y: -0.4688786
			z: 0.6559708
		}, Vertex{
			x: 0.1258684
			y: -0.4688786
			z: -0.6559708
		}]
		faces:     [[0, 36, 28, 48, 12], [1, 37, 29, 49, 13],
			[2, 38, 30, 50, 14], [3, 39, 31, 51, 15], [4, 40, 32, 53, 17],
			[5, 41, 33, 52, 16], [6, 42, 34, 55, 19], [7, 43, 35, 54, 18],
			[8, 44, 24, 58, 22], [9, 45, 25, 59, 23], [10, 46, 26, 56, 20],
			[11, 47, 27, 57, 21], [0, 2, 14], [1, 3, 15], [2, 0, 12],
			[3, 1, 13], [4, 5, 16], [5, 4, 17], [6, 7, 18], [7, 6, 19],
			[8, 11, 21], [9, 10, 20], [10, 9, 23], [11, 8, 22],
			[12, 48, 56], [13, 49, 57], [14, 50, 58], [15, 51, 59],
			[16, 52, 48], [17, 53, 49], [18, 54, 50], [19, 55, 51],
			[20, 56, 52], [21, 57, 53], [22, 58, 54], [23, 59, 55],
			[24, 44, 36], [25, 45, 37], [26, 46, 38], [27, 47, 39],
			[28, 36, 40], [29, 37, 41], [30, 38, 42], [31, 39, 43],
			[32, 40, 44], [33, 41, 45], [34, 42, 46], [35, 43, 47],
			[36, 0, 24], [37, 1, 25], [38, 2, 26], [39, 3, 27],
			[40, 4, 28], [41, 5, 29], [42, 6, 30], [43, 7, 31],
			[44, 8, 32], [45, 9, 33], [46, 10, 34], [47, 11, 35],
			[48, 28, 16], [49, 29, 17], [50, 30, 18], [51, 31, 19],
			[52, 33, 20], [53, 32, 21], [54, 35, 22], [55, 34, 23],
			[56, 26, 12], [57, 27, 13], [58, 24, 14], [59, 25, 15],
			[24, 0, 14], [25, 1, 15], [26, 2, 12], [27, 3, 13],
			[28, 4, 16], [29, 5, 17], [30, 6, 18], [31, 7, 19],
			[32, 8, 21], [33, 9, 20], [34, 10, 23], [35, 11, 22],
			[36, 44, 40], [37, 45, 41], [38, 46, 42], [39, 47, 43],
			[48, 52, 56], [49, 53, 57], [50, 54, 58], [51, 55, 59]]
	},
	Polyhedron{
		name:      'GreatIcosicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.1909830
			z: 1.118034
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: -1.118034
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: 1.118034
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: 1.118034
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: -1.118034
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: -1.118034
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: 0.1909830
			y: 1.118034
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: -1.118034
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: 1.118034
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: -1.118034
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: 1.0
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: -1.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: 1.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: -1.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: 1.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: -1.0
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: 1.0
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: 1.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: 1.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: 1.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: -1.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: -1.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: -1.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: -1.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: 1.0
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: -1.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: -1.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: 1.0
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: 1.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: -1.0
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: -1.0
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: 0.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: 0.618034
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: -0.618034
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: -0.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: 0.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: 0.618034
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: -0.618034
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: -0.618034
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: 0.618034
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: -0.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: 0.618034
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: -0.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: 0.618034
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: -0.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: 0.618034
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: 0.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: 0.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: 0.618034
			y: -0.809017
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: -0.618034
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: -0.618034
			y: -0.809017
			z: -0.5
		}]
		faces:     [[0, 42, 11, 55, 5, 44], [0, 48, 7, 59, 9, 38],
			[1, 39, 9, 58, 6, 49], [1, 45, 4, 54, 11, 43], [2, 36, 8, 57, 7, 50],
			[2, 46, 5, 53, 10, 40], [3, 41, 10, 52, 4, 47], [3, 51, 6, 56, 8, 37],
			[15, 13, 29, 44, 46, 31], [15, 23, 22, 14, 58, 59],
			[18, 16, 32, 49, 51, 34], [18, 26, 27, 19, 55, 54],
			[20, 21, 13, 57, 56, 12], [20, 28, 32, 24, 42, 38],
			[25, 24, 16, 52, 53, 17], [25, 33, 29, 21, 39, 43],
			[30, 22, 36, 40, 26, 34], [30, 47, 45, 28, 12, 14],
			[35, 27, 41, 37, 23, 31], [35, 50, 48, 33, 17, 19],
			[0, 44, 29, 33, 48], [1, 49, 32, 28, 45], [2, 50, 35, 31, 46],
			[3, 47, 30, 34, 51], [4, 52, 16, 18, 54], [5, 55, 19, 17, 53],
			[6, 58, 14, 12, 56], [7, 57, 13, 15, 59], [8, 36, 22, 23, 37],
			[9, 39, 21, 20, 38], [10, 41, 27, 26, 40], [11, 42, 24, 25, 43],
			[0, 38, 42], [1, 43, 39], [2, 40, 36], [3, 37, 41],
			[4, 45, 47], [5, 46, 44], [6, 51, 49], [7, 48, 50],
			[8, 56, 57], [9, 59, 58], [10, 53, 52], [11, 54, 55],
			[12, 28, 20], [13, 21, 29], [14, 22, 30], [15, 31, 23],
			[16, 24, 32], [17, 33, 25], [18, 34, 26], [19, 27, 35]]
	},
	Polyhedron{
		name:      'SmallRhombihexacron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 3.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -3.414214
		}, Vertex{
			x: 3.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -3.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 3.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -3.414214
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[0, 10, 2, 14], [0, 11, 5, 6], [0, 12, 4, 8],
			[0, 13, 3, 16], [1, 10, 4, 7], [1, 11, 2, 17], [1, 12, 3, 15],
			[1, 13, 5, 9], [2, 14, 4, 6], [2, 15, 1, 10], [2, 16, 0, 11],
			[2, 17, 5, 7], [3, 14, 0, 12], [3, 15, 4, 9], [3, 16, 5, 8],
			[3, 17, 1, 13], [4, 6, 0, 10], [4, 7, 2, 15], [4, 8, 3, 14],
			[4, 9, 1, 12], [5, 6, 2, 16], [5, 7, 1, 11], [5, 8, 0, 13],
			[5, 9, 3, 17]]
	},
	Polyhedron{
		name:      'SmallRhombidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 2.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -2.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 2.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -2.118034
		}, Vertex{
			x: 2.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 2.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 2.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -2.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -2.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 2.118034
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -2.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 2.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -2.118034
			z: -0.5
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: 1.618034
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: -1.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: 1.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: -1.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: 1.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: -1.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: 1.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: 1.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: 1.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: 1.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: -1.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: -1.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: -1.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: -1.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: 1.618034
			z: -1.309017
		}, Vertex{
			x: 0.809017
			y: -1.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: -1.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: 1.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: 1.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: -1.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: -1.618034
			z: -1.309017
		}]
		faces:     [[0, 24, 56, 48, 12, 14, 50, 58, 26, 2], [0, 36, 44, 32, 17, 21, 34, 48, 40,
			4],
			[7, 3, 39, 47, 33, 18, 22, 35, 51, 43], [7, 5, 25, 53, 45, 9, 11, 47, 55, 27],
			[10, 8, 44, 52, 24, 4, 6, 26, 54, 46], [10, 11, 29, 37, 53, 17, 16, 52, 36, 28],
			[13, 31, 43, 59, 23, 22, 58, 42, 30, 12], [13, 49, 57, 25, 1, 3, 27, 59, 51, 15],
			[19, 33, 46, 38, 2, 6, 42, 50, 35, 23], [19, 55, 39, 29, 9, 8, 28, 38, 54, 18],
			[20, 16, 32, 45, 37, 1, 5, 41, 49, 34], [20, 21, 57, 41, 31, 15, 14, 30, 40, 56],
			[24, 0, 36, 52], [24, 56, 40, 4], [25, 5, 41, 57],
			[25, 53, 37, 1], [26, 6, 42, 58], [26, 54, 38, 2],
			[27, 3, 39, 55], [27, 59, 43, 7], [28, 8, 44, 36],
			[28, 38, 46, 10], [29, 11, 47, 39], [29, 37, 45, 9],
			[30, 14, 50, 42], [30, 40, 48, 12], [31, 13, 49, 41],
			[31, 43, 51, 15], [32, 16, 52, 44], [32, 45, 53, 17],
			[33, 19, 55, 47], [33, 46, 54, 18], [34, 21, 57, 49],
			[34, 48, 56, 20], [35, 22, 58, 50], [35, 51, 59, 23],
			[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9], [12, 13, 15, 14],
			[16, 17, 21, 20], [18, 22, 23, 19]]
	},
	Polyhedron{
		name:      'GreatInvertedPentagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.1533576
			y: 0.3791678
			z: -0.4074937
		}, Vertex{
			x: -0.1533576
			y: 0.3791678
			z: 0.4074937
		}, Vertex{
			x: -0.1533576
			y: -0.3791678
			z: -0.4074937
		}, Vertex{
			x: 0.1533576
			y: -0.3791678
			z: 0.4074937
		}, Vertex{
			x: 0.3791678
			y: -0.4074937
			z: 0.1533576
		}, Vertex{
			x: -0.3791678
			y: -0.4074937
			z: -0.1533576
		}, Vertex{
			x: -0.3791678
			y: 0.4074937
			z: 0.1533576
		}, Vertex{
			x: 0.3791678
			y: 0.4074937
			z: -0.1533576
		}, Vertex{
			x: -0.4074937
			y: 0.1533576
			z: 0.3791678
		}, Vertex{
			x: 0.4074937
			y: 0.1533576
			z: -0.3791678
		}, Vertex{
			x: 0.4074937
			y: -0.1533576
			z: 0.3791678
		}, Vertex{
			x: -0.4074937
			y: -0.1533576
			z: -0.3791678
		}, Vertex{
			x: 0.5393484
			y: 0.0
			z: 0.2060127
		}, Vertex{
			x: 0.5393484
			y: 0.0
			z: -0.2060127
		}, Vertex{
			x: -0.5393484
			y: 0.0
			z: 0.2060127
		}, Vertex{
			x: -0.5393484
			y: 0.0
			z: -0.2060127
		}, Vertex{
			x: 0.0
			y: 0.2060127
			z: 0.5393484
		}, Vertex{
			x: 0.0
			y: 0.2060127
			z: -0.5393484
		}, Vertex{
			x: 0.0
			y: -0.2060127
			z: 0.5393484
		}, Vertex{
			x: 0.0
			y: -0.2060127
			z: -0.5393484
		}, Vertex{
			x: 0.2060127
			y: 0.5393484
			z: 0.0
		}, Vertex{
			x: -0.2060127
			y: 0.5393484
			z: 0.0
		}, Vertex{
			x: 0.2060127
			y: -0.5393484
			z: 0.0
		}, Vertex{
			x: -0.2060127
			y: -0.5393484
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.3779726
			z: -0.2335999
		}, Vertex{
			x: 0.0
			y: 0.3779726
			z: 0.2335999
		}, Vertex{
			x: 0.0
			y: -0.3779726
			z: -0.2335999
		}, Vertex{
			x: 0.0
			y: -0.3779726
			z: 0.2335999
		}, Vertex{
			x: 0.3779726
			y: -0.2335999
			z: 0.0
		}, Vertex{
			x: -0.3779726
			y: -0.2335999
			z: 0.0
		}, Vertex{
			x: 0.3779726
			y: 0.2335999
			z: 0.0
		}, Vertex{
			x: -0.3779726
			y: 0.2335999
			z: 0.0
		}, Vertex{
			x: -0.2335999
			y: 0.0
			z: 0.3779726
		}, Vertex{
			x: -0.2335999
			y: 0.0
			z: -0.3779726
		}, Vertex{
			x: 0.2335999
			y: 0.0
			z: 0.3779726
		}, Vertex{
			x: 0.2335999
			y: 0.0
			z: -0.3779726
		}, Vertex{
			x: -0.03749140
			y: 0.5666434
			z: -0.1041519
		}, Vertex{
			x: 0.03749140
			y: 0.5666434
			z: 0.1041519
		}, Vertex{
			x: 0.03749140
			y: -0.5666434
			z: -0.1041519
		}, Vertex{
			x: -0.03749140
			y: -0.5666434
			z: 0.1041519
		}, Vertex{
			x: -0.5666434
			y: -0.1041519
			z: 0.03749140
		}, Vertex{
			x: 0.5666434
			y: -0.1041519
			z: -0.03749140
		}, Vertex{
			x: 0.5666434
			y: 0.1041519
			z: 0.03749140
		}, Vertex{
			x: -0.5666434
			y: 0.1041519
			z: -0.03749140
		}, Vertex{
			x: 0.1041519
			y: 0.03749140
			z: 0.5666434
		}, Vertex{
			x: -0.1041519
			y: 0.03749140
			z: -0.5666434
		}, Vertex{
			x: -0.1041519
			y: -0.03749140
			z: 0.5666434
		}, Vertex{
			x: 0.1041519
			y: -0.03749140
			z: -0.5666434
		}, Vertex{
			x: -0.1968472
			y: 0.1874755
			z: 0.5093545
		}, Vertex{
			x: 0.1968472
			y: 0.1874755
			z: -0.5093545
		}, Vertex{
			x: 0.1968472
			y: -0.1874755
			z: 0.5093545
		}, Vertex{
			x: -0.1968472
			y: -0.1874755
			z: -0.5093545
		}, Vertex{
			x: 0.1874755
			y: 0.5093545
			z: -0.1968472
		}, Vertex{
			x: -0.1874755
			y: 0.5093545
			z: 0.1968472
		}, Vertex{
			x: -0.1874755
			y: -0.5093545
			z: -0.1968472
		}, Vertex{
			x: 0.1874755
			y: -0.5093545
			z: 0.1968472
		}, Vertex{
			x: 0.5093545
			y: -0.1968472
			z: 0.1874755
		}, Vertex{
			x: -0.5093545
			y: -0.1968472
			z: -0.1874755
		}, Vertex{
			x: -0.5093545
			y: 0.1968472
			z: 0.1874755
		}, Vertex{
			x: 0.5093545
			y: 0.1968472
			z: -0.1874755
		}, Vertex{
			x: -0.2106465
			y: 0.4718631
			z: -0.2575096
		}, Vertex{
			x: 0.2106465
			y: 0.4718631
			z: 0.2575096
		}, Vertex{
			x: 0.2106465
			y: -0.4718631
			z: -0.2575096
		}, Vertex{
			x: -0.2106465
			y: -0.4718631
			z: 0.2575096
		}, Vertex{
			x: 0.4718631
			y: -0.2575096
			z: -0.2106465
		}, Vertex{
			x: -0.4718631
			y: -0.2575096
			z: 0.2106465
		}, Vertex{
			x: -0.4718631
			y: 0.2575096
			z: -0.2106465
		}, Vertex{
			x: 0.4718631
			y: 0.2575096
			z: 0.2106465
		}, Vertex{
			x: -0.2575096
			y: -0.2106465
			z: 0.4718631
		}, Vertex{
			x: 0.2575096
			y: -0.2106465
			z: -0.4718631
		}, Vertex{
			x: 0.2575096
			y: 0.2106465
			z: 0.4718631
		}, Vertex{
			x: -0.2575096
			y: 0.2106465
			z: -0.4718631
		}, Vertex{
			x: 0.4449851
			y: 0.09269529
			z: 0.3559969
		}, Vertex{
			x: -0.4449851
			y: 0.09269529
			z: -0.3559969
		}, Vertex{
			x: -0.4449851
			y: -0.09269529
			z: 0.3559969
		}, Vertex{
			x: 0.4449851
			y: -0.09269529
			z: -0.3559969
		}, Vertex{
			x: -0.09269529
			y: 0.3559969
			z: -0.4449851
		}, Vertex{
			x: 0.09269529
			y: 0.3559969
			z: 0.4449851
		}, Vertex{
			x: 0.09269529
			y: -0.3559969
			z: -0.4449851
		}, Vertex{
			x: -0.09269529
			y: -0.3559969
			z: 0.4449851
		}, Vertex{
			x: -0.3559969
			y: -0.4449851
			z: 0.09269529
		}, Vertex{
			x: 0.3559969
			y: -0.4449851
			z: -0.09269529
		}, Vertex{
			x: 0.3559969
			y: 0.4449851
			z: 0.09269529
		}, Vertex{
			x: -0.3559969
			y: 0.4449851
			z: -0.09269529
		}, Vertex{
			x: -0.3333356
			y: -0.3333356
			z: -0.3333356
		}, Vertex{
			x: -0.3333356
			y: -0.3333356
			z: 0.3333356
		}, Vertex{
			x: 0.3333356
			y: -0.3333356
			z: -0.3333356
		}, Vertex{
			x: 0.3333356
			y: -0.3333356
			z: 0.3333356
		}, Vertex{
			x: -0.3333356
			y: 0.3333356
			z: -0.3333356
		}, Vertex{
			x: -0.3333356
			y: 0.3333356
			z: 0.3333356
		}, Vertex{
			x: 0.3333356
			y: 0.3333356
			z: -0.3333356
		}, Vertex{
			x: 0.3333356
			y: 0.3333356
			z: 0.3333356
		}]
		faces:     [[24, 0, 2, 14, 36], [24, 36, 72, 86, 76],
			[24, 76, 40, 16, 52], [24, 52, 64, 84, 60], [24, 60, 48, 12, 0],
			[25, 1, 3, 13, 37], [25, 37, 73, 85, 77], [25, 77, 41, 17, 53],
			[25, 53, 65, 87, 61], [25, 61, 49, 15, 1], [26, 2, 0, 12, 38],
			[26, 38, 74, 88, 78], [26, 78, 42, 18, 54], [26, 54, 66, 90, 62],
			[26, 62, 50, 14, 2], [27, 3, 1, 15, 39], [27, 39, 75, 91, 79],
			[27, 79, 43, 19, 55], [27, 55, 67, 89, 63], [27, 63, 51, 13, 3],
			[28, 4, 5, 17, 41], [28, 41, 77, 85, 81], [28, 81, 45, 20, 56],
			[28, 56, 68, 84, 64], [28, 64, 52, 16, 4], [29, 5, 4, 16, 40],
			[29, 40, 76, 86, 80], [29, 80, 44, 21, 57], [29, 57, 69, 87, 65],
			[29, 65, 53, 17, 5], [30, 7, 6, 18, 42], [30, 42, 78, 88, 82],
			[30, 82, 46, 22, 59], [30, 59, 71, 89, 67], [30, 67, 55, 19, 7],
			[31, 6, 7, 19, 43], [31, 43, 79, 91, 83], [31, 83, 47, 23, 58],
			[31, 58, 70, 90, 66], [31, 66, 54, 18, 6], [32, 8, 11, 22, 46],
			[32, 46, 82, 88, 74], [32, 74, 38, 12, 48], [32, 48, 60, 84, 68],
			[32, 68, 56, 20, 8], [33, 11, 8, 20, 45], [33, 45, 81, 85, 73],
			[33, 73, 37, 13, 51], [33, 51, 63, 89, 71], [33, 71, 59, 22, 11],
			[34, 10, 9, 21, 44], [34, 44, 80, 86, 72], [34, 72, 36, 14, 50],
			[34, 50, 62, 90, 70], [34, 70, 58, 23, 10], [35, 9, 10, 23, 47],
			[35, 47, 83, 91, 75], [35, 75, 39, 15, 49], [35, 49, 61, 87, 69],
			[35, 69, 57, 21, 9]]
	},
	Polyhedron{
		name:      'UniformGreatRhombicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -0.1909830
		}, Vertex{
			x: 0.690983
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: -0.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: 0.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: -0.618034
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.1909830
			y: -0.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: -0.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: -0.618034
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: -0.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: 0.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: 0.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.618034
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.618034
			z: 0.309017
		}, Vertex{
			x: -0.618034
			y: -0.309017
			z: 0.1909830
		}, Vertex{
			x: -0.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.618034
			y: -0.309017
			z: 0.1909830
		}, Vertex{
			x: 0.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: -0.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: -0.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: 0.618034
			y: 0.309017
			z: -0.1909830
		}]
		faces:     [[24, 52, 16, 20, 56], [25, 57, 21, 17, 53],
			[26, 58, 22, 18, 54], [27, 55, 19, 23, 59], [28, 36, 0, 2, 38],
			[29, 39, 3, 1, 37], [30, 42, 6, 4, 40], [31, 41, 5, 7, 43],
			[32, 44, 8, 9, 45], [33, 47, 11, 10, 46], [34, 49, 13, 12, 48],
			[35, 50, 14, 15, 51], [0, 36, 52, 24], [1, 25, 53, 37],
			[2, 26, 54, 38], [3, 39, 55, 27], [4, 24, 56, 40],
			[5, 41, 57, 25], [6, 42, 58, 26], [7, 27, 59, 43],
			[8, 44, 36, 28], [9, 29, 37, 45], [10, 28, 38, 46],
			[11, 47, 39, 29], [12, 30, 40, 48], [13, 49, 41, 31],
			[14, 50, 42, 30], [15, 31, 43, 51], [16, 52, 44, 32],
			[17, 32, 45, 53], [18, 33, 46, 54], [19, 55, 47, 33],
			[20, 34, 48, 56], [21, 57, 49, 34], [22, 58, 50, 35],
			[23, 35, 51, 59], [0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9],
			[12, 13, 15, 14], [16, 17, 21, 20], [18, 22, 23, 19],
			[24, 4, 0], [25, 1, 5], [26, 2, 6], [27, 7, 3], [28, 10, 8],
			[29, 9, 11], [30, 12, 14], [31, 15, 13], [32, 17, 16],
			[33, 18, 19], [34, 20, 21], [35, 23, 22], [36, 44, 52],
			[37, 53, 45], [38, 54, 46], [39, 47, 55], [40, 56, 48],
			[41, 49, 57], [42, 50, 58], [43, 59, 51]]
	},
	Polyhedron{
		name:      'SmallHexagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.309017
			y: 0.0
			z: 1.366760
		}, Vertex{
			x: 0.309017
			y: 0.0
			z: -1.366760
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: 1.366760
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: -1.366760
		}, Vertex{
			x: 1.366760
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: 1.366760
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: -1.366760
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: -1.366760
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.366760
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: 1.366760
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: -1.366760
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: -1.366760
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 0.5768607
			y: 0.4333802
			z: 1.201224
		}, Vertex{
			x: 0.5768607
			y: 0.4333802
			z: -1.201224
		}, Vertex{
			x: 0.5768607
			y: -0.4333802
			z: 1.201224
		}, Vertex{
			x: 0.5768607
			y: -0.4333802
			z: -1.201224
		}, Vertex{
			x: -0.5768607
			y: 0.4333802
			z: 1.201224
		}, Vertex{
			x: -0.5768607
			y: 0.4333802
			z: -1.201224
		}, Vertex{
			x: -0.5768607
			y: -0.4333802
			z: 1.201224
		}, Vertex{
			x: -0.5768607
			y: -0.4333802
			z: -1.201224
		}, Vertex{
			x: 1.201224
			y: 0.5768607
			z: 0.4333802
		}, Vertex{
			x: 1.201224
			y: 0.5768607
			z: -0.4333802
		}, Vertex{
			x: 1.201224
			y: -0.5768607
			z: 0.4333802
		}, Vertex{
			x: 1.201224
			y: -0.5768607
			z: -0.4333802
		}, Vertex{
			x: -1.201224
			y: 0.5768607
			z: 0.4333802
		}, Vertex{
			x: -1.201224
			y: 0.5768607
			z: -0.4333802
		}, Vertex{
			x: -1.201224
			y: -0.5768607
			z: 0.4333802
		}, Vertex{
			x: -1.201224
			y: -0.5768607
			z: -0.4333802
		}, Vertex{
			x: 0.4333802
			y: 1.201224
			z: 0.5768607
		}, Vertex{
			x: 0.4333802
			y: 1.201224
			z: -0.5768607
		}, Vertex{
			x: 0.4333802
			y: -1.201224
			z: 0.5768607
		}, Vertex{
			x: 0.4333802
			y: -1.201224
			z: -0.5768607
		}, Vertex{
			x: -0.4333802
			y: 1.201224
			z: 0.5768607
		}, Vertex{
			x: -0.4333802
			y: 1.201224
			z: -0.5768607
		}, Vertex{
			x: -0.4333802
			y: -1.201224
			z: 0.5768607
		}, Vertex{
			x: -0.4333802
			y: -1.201224
			z: -0.5768607
		}, Vertex{
			x: 0.7252591
			y: 0.0
			z: 1.173494
		}, Vertex{
			x: 0.7252591
			y: 0.0
			z: -1.173494
		}, Vertex{
			x: -0.7252591
			y: 0.0
			z: 1.173494
		}, Vertex{
			x: -0.7252591
			y: 0.0
			z: -1.173494
		}, Vertex{
			x: 1.173494
			y: 0.7252591
			z: 0.0
		}, Vertex{
			x: 1.173494
			y: -0.7252591
			z: 0.0
		}, Vertex{
			x: -1.173494
			y: 0.7252591
			z: 0.0
		}, Vertex{
			x: -1.173494
			y: -0.7252591
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.173494
			z: 0.7252591
		}, Vertex{
			x: 0.0
			y: 1.173494
			z: -0.7252591
		}, Vertex{
			x: 0.0
			y: -1.173494
			z: 0.7252591
		}, Vertex{
			x: 0.0
			y: -1.173494
			z: -0.7252591
		}, Vertex{
			x: 0.2678437
			y: 0.9333802
			z: 1.010241
		}, Vertex{
			x: 0.2678437
			y: 0.9333802
			z: -1.010241
		}, Vertex{
			x: 0.2678437
			y: -0.9333802
			z: 1.010241
		}, Vertex{
			x: 0.2678437
			y: -0.9333802
			z: -1.010241
		}, Vertex{
			x: -0.2678437
			y: 0.9333802
			z: 1.010241
		}, Vertex{
			x: -0.2678437
			y: 0.9333802
			z: -1.010241
		}, Vertex{
			x: -0.2678437
			y: -0.9333802
			z: 1.010241
		}, Vertex{
			x: -0.2678437
			y: -0.9333802
			z: -1.010241
		}, Vertex{
			x: 1.010241
			y: 0.2678437
			z: 0.9333802
		}, Vertex{
			x: 1.010241
			y: 0.2678437
			z: -0.9333802
		}, Vertex{
			x: 1.010241
			y: -0.2678437
			z: 0.9333802
		}, Vertex{
			x: 1.010241
			y: -0.2678437
			z: -0.9333802
		}, Vertex{
			x: -1.010241
			y: 0.2678437
			z: 0.9333802
		}, Vertex{
			x: -1.010241
			y: 0.2678437
			z: -0.9333802
		}, Vertex{
			x: -1.010241
			y: -0.2678437
			z: 0.9333802
		}, Vertex{
			x: -1.010241
			y: -0.2678437
			z: -0.9333802
		}, Vertex{
			x: 0.9333802
			y: 1.010241
			z: 0.2678437
		}, Vertex{
			x: 0.9333802
			y: 1.010241
			z: -0.2678437
		}, Vertex{
			x: 0.9333802
			y: -1.010241
			z: 0.2678437
		}, Vertex{
			x: 0.9333802
			y: -1.010241
			z: -0.2678437
		}, Vertex{
			x: -0.9333802
			y: 1.010241
			z: 0.2678437
		}, Vertex{
			x: -0.9333802
			y: 1.010241
			z: -0.2678437
		}, Vertex{
			x: -0.9333802
			y: -1.010241
			z: 0.2678437
		}, Vertex{
			x: -0.9333802
			y: -1.010241
			z: -0.2678437
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: -0.809017
		}]
		faces:     [[60, 0, 17, 74, 100, 82], [60, 82, 20, 44, 97, 36],
			[60, 36, 12, 2, 16, 38], [60, 38, 101, 46, 21, 80],
			[60, 80, 96, 72, 13, 0], [61, 1, 15, 73, 98, 81],
			[61, 81, 22, 47, 103, 39], [61, 39, 18, 3, 14, 37],
			[61, 37, 99, 45, 23, 83], [61, 83, 102, 75, 19, 1],
			[62, 2, 12, 76, 104, 84], [62, 84, 25, 50, 109, 42],
			[62, 42, 17, 0, 13, 40], [62, 40, 105, 48, 24, 86],
			[62, 86, 108, 78, 16, 2], [63, 3, 18, 79, 110, 87],
			[63, 87, 27, 49, 107, 41], [63, 41, 15, 1, 19, 43],
			[63, 43, 111, 51, 26, 85], [63, 85, 106, 77, 14, 3],
			[64, 4, 22, 81, 98, 89], [64, 89, 29, 52, 97, 44],
			[64, 44, 20, 5, 23, 45], [64, 45, 99, 53, 28, 88],
			[64, 88, 96, 80, 21, 4], [65, 5, 20, 82, 100, 90],
			[65, 90, 31, 55, 103, 47], [65, 47, 22, 4, 21, 46],
			[65, 46, 101, 54, 30, 91], [65, 91, 102, 83, 23, 5],
			[66, 6, 25, 84, 104, 92], [66, 92, 32, 57, 107, 49],
			[66, 49, 27, 7, 24, 48], [66, 48, 105, 56, 33, 93],
			[66, 93, 106, 85, 26, 6], [67, 7, 27, 87, 110, 95],
			[67, 95, 34, 58, 109, 50], [67, 50, 25, 6, 26, 51],
			[67, 51, 111, 59, 35, 94], [67, 94, 108, 86, 24, 7],
			[68, 8, 32, 92, 104, 76], [68, 76, 12, 36, 97, 52],
			[68, 52, 29, 9, 33, 56], [68, 56, 105, 40, 13, 72],
			[68, 72, 96, 88, 28, 8], [69, 9, 29, 89, 98, 73],
			[69, 73, 15, 41, 107, 57], [69, 57, 32, 8, 28, 53],
			[69, 53, 99, 37, 14, 77], [69, 77, 106, 93, 33, 9],
			[70, 10, 31, 90, 100, 74], [70, 74, 17, 42, 109, 58],
			[70, 58, 34, 11, 30, 54], [70, 54, 101, 38, 16, 78],
			[70, 78, 108, 94, 35, 10], [71, 11, 34, 95, 110, 79],
			[71, 79, 18, 39, 103, 55], [71, 55, 31, 10, 35, 59],
			[71, 59, 111, 43, 19, 75], [71, 75, 102, 91, 30, 11]]
	},
	Polyhedron{
		name:      'MedialRhombicTriacontahedron'
		vertexes_: [Vertex{
			x: 0.75
			y: 0.0
			z: 1.213526
		}, Vertex{
			x: 0.75
			y: 0.0
			z: -1.213526
		}, Vertex{
			x: -0.75
			y: 0.0
			z: 1.213526
		}, Vertex{
			x: -0.75
			y: 0.0
			z: -1.213526
		}, Vertex{
			x: 1.213526
			y: 0.75
			z: 0.0
		}, Vertex{
			x: 1.213526
			y: -0.75
			z: 0.0
		}, Vertex{
			x: -1.213526
			y: 0.75
			z: 0.0
		}, Vertex{
			x: -1.213526
			y: -0.75
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.213526
			z: 0.75
		}, Vertex{
			x: 0.0
			y: 1.213526
			z: -0.75
		}, Vertex{
			x: 0.0
			y: -1.213526
			z: 0.75
		}, Vertex{
			x: 0.0
			y: -1.213526
			z: -0.75
		}, Vertex{
			x: 0.4635255
			y: 0.0
			z: 0.75
		}, Vertex{
			x: 0.4635255
			y: 0.0
			z: -0.75
		}, Vertex{
			x: -0.4635255
			y: 0.0
			z: 0.75
		}, Vertex{
			x: -0.4635255
			y: 0.0
			z: -0.75
		}, Vertex{
			x: 0.75
			y: 0.4635255
			z: 0.0
		}, Vertex{
			x: 0.75
			y: -0.4635255
			z: 0.0
		}, Vertex{
			x: -0.75
			y: 0.4635255
			z: 0.0
		}, Vertex{
			x: -0.75
			y: -0.4635255
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.75
			z: 0.4635255
		}, Vertex{
			x: 0.0
			y: 0.75
			z: -0.4635255
		}, Vertex{
			x: 0.0
			y: -0.75
			z: 0.4635255
		}, Vertex{
			x: 0.0
			y: -0.75
			z: -0.4635255
		}]
		faces:     [[0, 14, 7, 22], [0, 22, 11, 17], [0, 17, 1, 16],
			[0, 16, 9, 20], [0, 20, 6, 14], [3, 13, 5, 23], [3, 23, 10, 19],
			[3, 19, 2, 18], [3, 18, 8, 21], [3, 21, 4, 13], [1, 15, 6, 21],
			[1, 21, 8, 16], [2, 19, 11, 22], [2, 22, 5, 12], [4, 21, 6, 20],
			[4, 20, 2, 12], [5, 13, 9, 16], [5, 16, 8, 12], [6, 15, 11, 19],
			[6, 19, 10, 14], [7, 15, 1, 23], [7, 23, 5, 22], [8, 18, 7, 14],
			[8, 14, 10, 12], [9, 15, 7, 18], [9, 18, 2, 20], [10, 23, 1, 17],
			[10, 17, 4, 12], [11, 15, 9, 13], [11, 13, 4, 17]]
	},
	Polyhedron{
		name:      'SmallCubicuboctahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: -0.5
		}]
		faces:     [[0, 2, 18, 19, 3, 1, 17, 16], [0, 8, 9, 1, 5, 13, 12, 4],
			[11, 10, 2, 6, 14, 15, 7, 3], [11, 19, 23, 15, 13, 21, 17, 9],
			[20, 12, 14, 22, 18, 10, 8, 16], [20, 21, 5, 7, 23, 22, 6, 4],
			[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9], [12, 13, 15, 14],
			[16, 17, 21, 20], [18, 22, 23, 19], [0, 16, 8], [1, 9, 17],
			[2, 10, 18], [3, 19, 11], [4, 12, 20], [5, 21, 13],
			[6, 22, 14], [7, 15, 23]]
	},
	Polyhedron{
		name:      'SmallDodecicosahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.309017
			z: 1.618034
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: -1.618034
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: 1.618034
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: -1.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: 1.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: -1.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: 1.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: 1.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: 1.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 1.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: -1.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: -1.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: -1.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: -1.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: 1.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: 1.618034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: -1.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: -1.618034
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: 1.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: 1.618034
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: -1.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: -1.618034
			z: -0.5
		}, Vertex{
			x: 0.0
			y: 1.118034
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 1.118034
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -1.118034
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -1.118034
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 1.118034
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -1.118034
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 1.118034
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 1.118034
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 1.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 1.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 1.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: -1.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: -1.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: -1.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: -1.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 1.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 1.0
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: -1.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: -1.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 1.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 1.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: -1.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: -1.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 1.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: -1.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 1.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: -1.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 1.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: -1.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 1.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: -1.0
		}]
		faces:     [[0, 4, 30, 14, 51, 59, 55, 47, 10, 28], [0, 38, 46, 47, 39, 1, 25, 21, 20, 24],
			[2, 26, 22, 23, 27, 3, 37, 45, 44, 36], [2, 28, 8, 45, 53, 57, 49, 12, 30, 6],
			[5, 1, 29, 11, 46, 54, 58, 50, 15, 31], [5, 43, 51, 50, 42, 4, 24, 16, 17, 25],
			[7, 27, 19, 18, 26, 6, 40, 48, 49, 41], [7, 31, 13, 48, 56, 52, 44, 9, 29, 3],
			[33, 11, 9, 32, 16, 56, 40, 42, 58, 18], [33, 19, 59, 43, 41, 57, 17, 32, 8, 10],
			[34, 13, 15, 35, 22, 54, 38, 36, 52, 20], [34, 21, 53, 37, 39, 55, 23, 35, 14, 12],
			[0, 4, 42, 58, 54, 38], [0, 28, 8, 32, 16, 24], [3, 7, 41, 57, 53, 37],
			[3, 29, 11, 33, 19, 27], [17, 32, 9, 29, 1, 25], [17, 57, 49, 48, 56, 16],
			[18, 33, 10, 28, 2, 26], [18, 58, 50, 51, 59, 19],
			[34, 12, 30, 4, 24, 20], [34, 21, 25, 5, 31, 13],
			[35, 15, 31, 7, 27, 23], [35, 22, 26, 6, 30, 14],
			[40, 6, 2, 36, 52, 56], [40, 48, 13, 15, 50, 42],
			[43, 5, 1, 39, 55, 59], [43, 51, 14, 12, 49, 41],
			[44, 36, 38, 46, 11, 9], [44, 45, 53, 21, 20, 52],
			[47, 39, 37, 45, 8, 10], [47, 46, 54, 22, 23, 55]]
	},
	Polyhedron{
		name:      'SmallIcosicosidodecahedron'
		vertexes_: [Vertex{
			x: 1.309017
			y: 0.0
			z: -1.118034
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 1.118034
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -1.118034
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 1.118034
		}, Vertex{
			x: 0.0
			y: -1.118034
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -1.118034
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: 1.118034
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 1.118034
			z: -1.309017
		}, Vertex{
			x: -1.118034
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 1.118034
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -1.118034
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 1.118034
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 1.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: -1.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 1.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: -1.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 1.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: -1.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 1.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: -1.0
		}, Vertex{
			x: 1.309017
			y: 1.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 1.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 1.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 1.0
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: -1.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: -1.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: -1.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: -1.0
			z: -0.5
		}, Vertex{
			x: 1.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 1.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: -1.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: -1.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 1.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 1.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: -1.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: -1.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: -1.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: -1.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: 1.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: 1.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: -1.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: -1.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 1.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: 1.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: -1.618034
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: 1.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: -1.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: 1.618034
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: -1.618034
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: 1.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: -1.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: 1.618034
		}, Vertex{
			x: -0.309017
			y: -1.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: -1.618034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: -1.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: -1.618034
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: 1.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: 1.618034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 1.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: 1.618034
			z: -0.5
		}]
		faces:     [[0, 42, 11, 55, 5, 44], [0, 48, 7, 59, 9, 38],
			[1, 39, 9, 58, 6, 49], [1, 45, 4, 54, 11, 43], [2, 36, 8, 57, 7, 50],
			[2, 46, 5, 53, 10, 40], [3, 41, 10, 52, 4, 47], [3, 51, 6, 56, 8, 37],
			[15, 13, 29, 44, 46, 31], [15, 23, 22, 14, 58, 59],
			[18, 16, 32, 49, 51, 34], [18, 26, 27, 19, 55, 54],
			[20, 21, 13, 57, 56, 12], [20, 28, 32, 24, 42, 38],
			[25, 24, 16, 52, 53, 17], [25, 33, 29, 21, 39, 43],
			[30, 22, 36, 40, 26, 34], [30, 47, 45, 28, 12, 14],
			[35, 27, 41, 37, 23, 31], [35, 50, 48, 33, 17, 19],
			[0, 44, 29, 33, 48], [1, 49, 32, 28, 45], [2, 50, 35, 31, 46],
			[3, 47, 30, 34, 51], [4, 52, 16, 18, 54], [5, 55, 19, 17, 53],
			[6, 58, 14, 12, 56], [7, 57, 13, 15, 59], [8, 36, 22, 23, 37],
			[9, 39, 21, 20, 38], [10, 41, 27, 26, 40], [11, 42, 24, 25, 43],
			[0, 38, 42], [1, 43, 39], [2, 40, 36], [3, 37, 41],
			[4, 45, 47], [5, 46, 44], [6, 51, 49], [7, 48, 50],
			[8, 56, 57], [9, 59, 58], [10, 53, 52], [11, 54, 55],
			[12, 28, 20], [13, 21, 29], [14, 22, 30], [15, 31, 23],
			[16, 24, 32], [17, 33, 25], [18, 34, 26], [19, 27, 35]]
	},
	Polyhedron{
		name:      'DeltoidalIcositetrahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.414214
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: 0.7734591
			y: 0.7734591
			z: 0.7734591
		}, Vertex{
			x: 0.7734591
			y: 0.7734591
			z: -0.7734591
		}, Vertex{
			x: 0.7734591
			y: -0.7734591
			z: 0.7734591
		}, Vertex{
			x: 0.7734591
			y: -0.7734591
			z: -0.7734591
		}, Vertex{
			x: -0.7734591
			y: 0.7734591
			z: 0.7734591
		}, Vertex{
			x: -0.7734591
			y: 0.7734591
			z: -0.7734591
		}, Vertex{
			x: -0.7734591
			y: -0.7734591
			z: 0.7734591
		}, Vertex{
			x: -0.7734591
			y: -0.7734591
			z: -0.7734591
		}]
		faces:     [[0, 6, 18, 14], [0, 14, 22, 8], [0, 8, 24, 16],
			[0, 16, 20, 6], [1, 9, 23, 15], [1, 15, 19, 7], [1, 7, 21, 17],
			[1, 17, 25, 9], [2, 7, 19, 10], [2, 10, 18, 6], [2, 6, 20, 11],
			[2, 11, 21, 7], [3, 8, 22, 12], [3, 12, 23, 9], [3, 9, 25, 13],
			[3, 13, 24, 8], [4, 10, 19, 15], [4, 15, 23, 12],
			[4, 12, 22, 14], [4, 14, 18, 10], [5, 11, 20, 16],
			[5, 16, 24, 13], [5, 13, 25, 17], [5, 17, 21, 11]]
	},
	Polyhedron{
		name:      'TriakisTetrahedron'
		vertexes_: [Vertex{
			x: 1.060660
			y: 1.060660
			z: 1.060660
		}, Vertex{
			x: 1.060660
			y: -1.060660
			z: -1.060660
		}, Vertex{
			x: -1.060660
			y: -1.060660
			z: 1.060660
		}, Vertex{
			x: -1.060660
			y: 1.060660
			z: -1.060660
		}, Vertex{
			x: 0.6363961
			y: -0.6363961
			z: 0.6363961
		}, Vertex{
			x: 0.6363961
			y: 0.6363961
			z: -0.6363961
		}, Vertex{
			x: -0.6363961
			y: 0.6363961
			z: 0.6363961
		}, Vertex{
			x: -0.6363961
			y: -0.6363961
			z: -0.6363961
		}]
		faces:     [[4, 0, 2], [4, 2, 1], [4, 1, 0], [5, 0, 1],
			[5, 1, 3], [5, 3, 0], [6, 0, 3], [6, 3, 2], [6, 2, 0],
			[7, 1, 2], [7, 2, 3], [7, 3, 1]]
	},
	Polyhedron{
		name:      'CubitruncatedCuboctahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.2071068
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: 0.2071068
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 1.207107
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: -0.2071068
		}]
		faces:     [[0, 4, 26, 24, 6, 2, 28, 30], [1, 31, 29, 3, 7, 25, 27, 5],
			[8, 10, 33, 32, 11, 9, 34, 35], [12, 39, 38, 13, 15, 36, 37, 14],
			[16, 17, 44, 40, 21, 20, 41, 45], [18, 47, 43, 22, 23, 42, 46, 19],
			[0, 32, 33, 1, 5, 37, 36, 4], [2, 6, 38, 39, 7, 3, 35, 34],
			[8, 40, 44, 12, 14, 46, 42, 10], [9, 11, 43, 47, 15, 13, 45, 41],
			[16, 24, 26, 18, 19, 27, 25, 17], [20, 21, 29, 31, 23, 22, 30, 28],
			[0, 30, 22, 43, 11, 32], [1, 33, 10, 42, 23, 31],
			[2, 34, 9, 41, 20, 28], [3, 29, 21, 40, 8, 35], [4, 36, 15, 47, 18, 26],
			[5, 27, 19, 46, 14, 37], [6, 24, 16, 45, 13, 38],
			[7, 39, 12, 44, 17, 25]]
	},
	Polyhedron{
		name:      'MedialIcosacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.7783914
			y: 0.0
			z: 1.259464
		}, Vertex{
			x: 0.7783914
			y: 0.0
			z: -1.259464
		}, Vertex{
			x: -0.7783914
			y: 0.0
			z: 1.259464
		}, Vertex{
			x: -0.7783914
			y: 0.0
			z: -1.259464
		}, Vertex{
			x: 1.259464
			y: 0.7783914
			z: 0.0
		}, Vertex{
			x: 1.259464
			y: -0.7783914
			z: 0.0
		}, Vertex{
			x: -1.259464
			y: 0.7783914
			z: 0.0
		}, Vertex{
			x: -1.259464
			y: -0.7783914
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.259464
			z: 0.7783914
		}, Vertex{
			x: 0.0
			y: 1.259464
			z: -0.7783914
		}, Vertex{
			x: 0.0
			y: -1.259464
			z: 0.7783914
		}, Vertex{
			x: 0.0
			y: -1.259464
			z: -0.7783914
		}, Vertex{
			x: 0.6496271
			y: 0.0
			z: 1.051119
		}, Vertex{
			x: 0.6496271
			y: 0.0
			z: -1.051119
		}, Vertex{
			x: -0.6496271
			y: 0.0
			z: 1.051119
		}, Vertex{
			x: -0.6496271
			y: 0.0
			z: -1.051119
		}, Vertex{
			x: 1.051119
			y: 0.6496271
			z: 0.0
		}, Vertex{
			x: 1.051119
			y: -0.6496271
			z: 0.0
		}, Vertex{
			x: -1.051119
			y: 0.6496271
			z: 0.0
		}, Vertex{
			x: -1.051119
			y: -0.6496271
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.051119
			z: 0.6496271
		}, Vertex{
			x: 0.0
			y: 1.051119
			z: -0.6496271
		}, Vertex{
			x: 0.0
			y: -1.051119
			z: 0.6496271
		}, Vertex{
			x: 0.0
			y: -1.051119
			z: -0.6496271
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[12, 5, 28, 8], [12, 8, 32, 40], [12, 40, 26, 42],
			[12, 42, 34, 9], [12, 9, 29, 5], [13, 4, 29, 9], [13, 9, 35, 43],
			[13, 43, 27, 41], [13, 41, 33, 8], [13, 8, 28, 4],
			[14, 7, 31, 11], [14, 11, 34, 38], [14, 38, 24, 36],
			[14, 36, 32, 10], [14, 10, 30, 7], [15, 6, 30, 10],
			[15, 10, 33, 37], [15, 37, 25, 39], [15, 39, 35, 11],
			[15, 11, 31, 6], [16, 1, 33, 10], [16, 10, 32, 0],
			[16, 0, 24, 38], [16, 38, 29, 39], [16, 39, 25, 1],
			[17, 2, 34, 11], [17, 11, 35, 3], [17, 3, 25, 37],
			[17, 37, 28, 36], [17, 36, 24, 2], [18, 0, 32, 8],
			[18, 8, 33, 1], [18, 1, 27, 43], [18, 43, 31, 42],
			[18, 42, 26, 0], [19, 2, 26, 40], [19, 40, 30, 41],
			[19, 41, 27, 3], [19, 3, 35, 9], [19, 9, 34, 2], [20, 2, 24, 4],
			[20, 4, 28, 37], [20, 37, 33, 41], [20, 41, 30, 6],
			[20, 6, 26, 2], [21, 3, 27, 7], [21, 7, 30, 40], [21, 40, 32, 36],
			[21, 36, 28, 5], [21, 5, 25, 3], [22, 0, 26, 6], [22, 6, 31, 43],
			[22, 43, 35, 39], [22, 39, 29, 4], [22, 4, 24, 0],
			[23, 1, 25, 5], [23, 5, 29, 38], [23, 38, 34, 42],
			[23, 42, 31, 7], [23, 7, 27, 1]]
	},
	Polyhedron{
		name:      'SmallDitrigonalIcosidodecahedron'
		vertexes_: [Vertex{
			x: -0.809017
			y: 0.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: 0.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: 0.0
			z: -0.309017
		}, Vertex{
			x: 0.809017
			y: 0.0
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: 0.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: 0.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: 0.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.5
		}]
		faces:     [[0, 6, 19, 15, 4], [0, 8, 1, 19, 18], [0, 14, 15, 1, 10],
			[7, 1, 5, 14, 18], [7, 11, 14, 12, 10], [7, 16, 12, 5, 3],
			[9, 2, 16, 17, 3], [9, 5, 8, 16, 18], [9, 19, 17, 8, 4],
			[13, 12, 2, 11, 3], [13, 15, 11, 6, 10], [13, 17, 6, 2, 4],
			[0, 4, 8], [0, 10, 6], [0, 18, 14], [1, 7, 10], [1, 8, 5],
			[1, 15, 19], [2, 6, 11], [2, 9, 4], [2, 12, 16], [3, 5, 9],
			[3, 11, 7], [3, 17, 13], [4, 15, 13], [5, 12, 14],
			[6, 17, 19], [7, 18, 16], [8, 17, 16], [9, 18, 19],
			[10, 12, 13], [11, 15, 14]]
	},
	Polyhedron{
		name:      'TruncatedCuboctahedron'
		vertexes_: [Vertex{
			x: 1.207107
			y: 0.5
			z: 1.914214
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: -1.914214
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: 1.914214
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: -1.914214
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: 1.914214
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: -1.914214
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: 1.914214
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: -1.914214
		}, Vertex{
			x: 1.914214
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: 1.914214
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: 1.914214
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: 1.914214
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: -1.914214
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: -1.914214
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: -1.914214
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: -1.914214
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.914214
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: 1.914214
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: -1.914214
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: -1.914214
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: 1.914214
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: 1.914214
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: -1.914214
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: -1.914214
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: 1.914214
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: -1.914214
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: 1.914214
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: -1.914214
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: 1.914214
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: -1.914214
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: 1.914214
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: -1.914214
		}, Vertex{
			x: 1.914214
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: 1.914214
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: 1.914214
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: 1.914214
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: -1.914214
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: -1.914214
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: -1.914214
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: -1.914214
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 1.914214
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: 1.914214
			z: -0.5
		}, Vertex{
			x: 1.207107
			y: -1.914214
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: -1.914214
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: 1.914214
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: 1.914214
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: -1.914214
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: -1.914214
			z: -0.5
		}]
		faces:     [[0, 24, 28, 4, 6, 30, 26, 2], [1, 3, 27, 31, 7, 5, 29, 25],
			[8, 32, 34, 10, 11, 35, 33, 9], [12, 13, 37, 39, 15, 14, 38, 36],
			[16, 40, 41, 17, 21, 45, 44, 20], [18, 22, 46, 47, 23, 19, 43, 42],
			[0, 32, 8, 40, 16, 24], [1, 25, 17, 41, 9, 33], [2, 26, 18, 42, 10, 34],
			[3, 35, 11, 43, 19, 27], [4, 28, 20, 44, 12, 36],
			[5, 37, 13, 45, 21, 29], [6, 38, 14, 46, 22, 30],
			[7, 31, 23, 47, 15, 39], [0, 2, 34, 32], [1, 33, 35, 3],
			[4, 36, 38, 6], [5, 7, 39, 37], [8, 9, 41, 40], [10, 42, 43, 11],
			[12, 44, 45, 13], [14, 15, 47, 46], [16, 20, 28, 24],
			[17, 25, 29, 21], [18, 26, 30, 22], [19, 23, 31, 27]]
	},
	Polyhedron{
		name:      'GreatRhombihexacron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.5857865
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.5857865
		}, Vertex{
			x: 0.5857865
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.5857865
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.5857865
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.5857865
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[0, 10, 2, 14], [0, 11, 5, 6], [0, 12, 4, 8],
			[0, 13, 3, 16], [1, 10, 4, 7], [1, 11, 2, 17], [1, 12, 3, 15],
			[1, 13, 5, 9], [2, 14, 4, 6], [2, 15, 1, 10], [2, 16, 0, 11],
			[2, 17, 5, 7], [3, 14, 0, 12], [3, 15, 4, 9], [3, 16, 5, 8],
			[3, 17, 1, 13], [4, 6, 0, 10], [4, 7, 2, 15], [4, 8, 3, 14],
			[4, 9, 1, 12], [5, 6, 2, 16], [5, 7, 1, 11], [5, 8, 0, 13],
			[5, 9, 3, 17]]
	},
	Polyhedron{
		name:      'GreatDirhombicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.1817730
			y: 0.1429011
			z: 0.6682349
		}, Vertex{
			x: 0.1817730
			y: 0.1429011
			z: -0.6682349
		}, Vertex{
			x: 0.1817730
			y: -0.1429011
			z: 0.6682349
		}, Vertex{
			x: 0.1817730
			y: -0.1429011
			z: -0.6682349
		}, Vertex{
			x: -0.1817730
			y: 0.1429011
			z: 0.6682349
		}, Vertex{
			x: -0.1817730
			y: 0.1429011
			z: -0.6682349
		}, Vertex{
			x: -0.1817730
			y: -0.1429011
			z: 0.6682349
		}, Vertex{
			x: -0.1817730
			y: -0.1429011
			z: -0.6682349
		}, Vertex{
			x: 0.6682349
			y: 0.1817730
			z: 0.1429011
		}, Vertex{
			x: 0.6682349
			y: 0.1817730
			z: -0.1429011
		}, Vertex{
			x: 0.6682349
			y: -0.1817730
			z: 0.1429011
		}, Vertex{
			x: 0.6682349
			y: -0.1817730
			z: -0.1429011
		}, Vertex{
			x: -0.6682349
			y: 0.1817730
			z: 0.1429011
		}, Vertex{
			x: -0.6682349
			y: 0.1817730
			z: -0.1429011
		}, Vertex{
			x: -0.6682349
			y: -0.1817730
			z: 0.1429011
		}, Vertex{
			x: -0.6682349
			y: -0.1817730
			z: -0.1429011
		}, Vertex{
			x: 0.1429011
			y: 0.6682349
			z: 0.1817730
		}, Vertex{
			x: 0.1429011
			y: 0.6682349
			z: -0.1817730
		}, Vertex{
			x: 0.1429011
			y: -0.6682349
			z: 0.1817730
		}, Vertex{
			x: 0.1429011
			y: -0.6682349
			z: -0.1817730
		}, Vertex{
			x: -0.1429011
			y: 0.6682349
			z: 0.1817730
		}, Vertex{
			x: -0.1429011
			y: 0.6682349
			z: -0.1817730
		}, Vertex{
			x: -0.1429011
			y: -0.6682349
			z: 0.1817730
		}, Vertex{
			x: -0.1429011
			y: -0.6682349
			z: -0.1817730
		}, Vertex{
			x: 0.0
			y: 0.437016
			z: 0.5558929
		}, Vertex{
			x: 0.0
			y: 0.437016
			z: -0.5558929
		}, Vertex{
			x: 0.0
			y: -0.437016
			z: 0.5558929
		}, Vertex{
			x: 0.0
			y: -0.437016
			z: -0.5558929
		}, Vertex{
			x: 0.5558929
			y: 0.0
			z: 0.437016
		}, Vertex{
			x: 0.5558929
			y: 0.0
			z: -0.437016
		}, Vertex{
			x: -0.5558929
			y: 0.0
			z: 0.437016
		}, Vertex{
			x: -0.5558929
			y: 0.0
			z: -0.437016
		}, Vertex{
			x: 0.437016
			y: 0.5558929
			z: 0.0
		}, Vertex{
			x: 0.437016
			y: -0.5558929
			z: 0.0
		}, Vertex{
			x: -0.437016
			y: 0.5558929
			z: 0.0
		}, Vertex{
			x: -0.437016
			y: -0.5558929
			z: 0.0
		}, Vertex{
			x: 0.4129919
			y: 0.2312188
			z: 0.5253338
		}, Vertex{
			x: 0.4129919
			y: 0.2312188
			z: -0.5253338
		}, Vertex{
			x: 0.4129919
			y: -0.2312188
			z: 0.5253338
		}, Vertex{
			x: 0.4129919
			y: -0.2312188
			z: -0.5253338
		}, Vertex{
			x: -0.4129919
			y: 0.2312188
			z: 0.5253338
		}, Vertex{
			x: -0.4129919
			y: 0.2312188
			z: -0.5253338
		}, Vertex{
			x: -0.4129919
			y: -0.2312188
			z: 0.5253338
		}, Vertex{
			x: -0.4129919
			y: -0.2312188
			z: -0.5253338
		}, Vertex{
			x: 0.5253338
			y: 0.4129919
			z: 0.2312188
		}, Vertex{
			x: 0.5253338
			y: 0.4129919
			z: -0.2312188
		}, Vertex{
			x: 0.5253338
			y: -0.4129919
			z: 0.2312188
		}, Vertex{
			x: 0.5253338
			y: -0.4129919
			z: -0.2312188
		}, Vertex{
			x: -0.5253338
			y: 0.4129919
			z: 0.2312188
		}, Vertex{
			x: -0.5253338
			y: 0.4129919
			z: -0.2312188
		}, Vertex{
			x: -0.5253338
			y: -0.4129919
			z: 0.2312188
		}, Vertex{
			x: -0.5253338
			y: -0.4129919
			z: -0.2312188
		}, Vertex{
			x: 0.2312188
			y: 0.5253338
			z: 0.4129919
		}, Vertex{
			x: 0.2312188
			y: 0.5253338
			z: -0.4129919
		}, Vertex{
			x: 0.2312188
			y: -0.5253338
			z: 0.4129919
		}, Vertex{
			x: 0.2312188
			y: -0.5253338
			z: -0.4129919
		}, Vertex{
			x: -0.2312188
			y: 0.5253338
			z: 0.4129919
		}, Vertex{
			x: -0.2312188
			y: 0.5253338
			z: -0.4129919
		}, Vertex{
			x: -0.2312188
			y: -0.5253338
			z: 0.4129919
		}, Vertex{
			x: -0.2312188
			y: -0.5253338
			z: -0.4129919
		}]
		faces:     [[16, 10, 53, 36, 29], [16, 41, 45, 34, 1],
			[17, 11, 52, 37, 28], [17, 40, 44, 34, 0], [18, 8, 55, 38, 29],
			[18, 43, 47, 35, 3], [19, 9, 54, 39, 28], [19, 42, 46, 35, 2],
			[20, 14, 57, 40, 31], [20, 37, 49, 32, 5], [21, 15, 56, 41, 30],
			[21, 36, 48, 32, 4], [22, 12, 59, 42, 31], [22, 39, 51, 33, 7],
			[23, 13, 58, 43, 30], [23, 38, 50, 33, 6], [24, 10, 6, 44, 54],
			[24, 14, 2, 48, 58], [25, 11, 7, 45, 55], [25, 15, 3, 49, 59],
			[26, 8, 4, 46, 52], [26, 12, 0, 50, 56], [27, 9, 5, 47, 53],
			[27, 13, 1, 51, 57], [0, 12, 7, 11], [0, 34, 7, 33],
			[2, 14, 5, 9], [2, 35, 5, 32], [4, 8, 3, 15], [4, 32, 3, 35],
			[6, 10, 1, 13], [6, 33, 1, 34], [8, 18, 15, 21], [8, 26, 15, 25],
			[10, 16, 13, 23], [10, 24, 13, 27], [12, 22, 11, 17],
			[12, 26, 11, 25], [14, 20, 9, 19], [14, 24, 9, 27],
			[16, 1, 23, 6], [16, 29, 23, 30], [18, 3, 21, 4],
			[18, 29, 21, 30], [20, 5, 19, 2], [20, 31, 19, 28],
			[22, 7, 17, 0], [22, 31, 17, 28], [24, 54, 27, 57],
			[24, 58, 27, 53], [26, 52, 25, 59], [26, 56, 25, 55],
			[28, 37, 31, 42], [28, 39, 31, 40], [30, 41, 29, 38],
			[30, 43, 29, 36], [32, 48, 35, 47], [32, 49, 35, 46],
			[34, 44, 33, 51], [34, 45, 33, 50], [36, 21, 43, 18],
			[36, 47, 43, 48], [38, 23, 41, 16], [38, 45, 41, 50],
			[40, 17, 39, 22], [40, 51, 39, 44], [42, 19, 37, 20],
			[42, 49, 37, 46], [44, 6, 51, 1], [44, 57, 51, 54],
			[46, 4, 49, 3], [46, 59, 49, 52], [48, 2, 47, 5],
			[48, 53, 47, 58], [50, 0, 45, 7], [50, 55, 45, 56],
			[52, 11, 59, 12], [52, 42, 59, 37], [54, 9, 57, 14],
			[54, 40, 57, 39], [56, 15, 55, 8], [56, 38, 55, 41],
			[58, 13, 53, 10], [58, 36, 53, 43], [0, 11, 22], [0, 33, 45],
			[1, 10, 23], [1, 33, 44], [2, 9, 20], [2, 32, 47],
			[3, 8, 21], [3, 32, 46], [4, 15, 18], [4, 35, 49],
			[5, 14, 19], [5, 35, 48], [6, 13, 16], [6, 34, 51],
			[7, 12, 17], [7, 34, 50], [24, 53, 13], [24, 57, 9],
			[25, 52, 12], [25, 56, 8], [26, 55, 15], [26, 59, 11],
			[27, 54, 14], [27, 58, 10], [36, 18, 30], [36, 58, 47],
			[37, 19, 31], [37, 59, 46], [38, 16, 30], [38, 56, 45],
			[39, 17, 31], [39, 57, 44], [40, 22, 28], [40, 54, 51],
			[41, 23, 29], [41, 55, 50], [42, 20, 28], [42, 52, 49],
			[43, 21, 29], [43, 53, 48]]
	},
	Polyhedron{
		name:      'GreatDodecahemicosahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: -0.309017
		}]
		faces:     [[0, 14, 15, 1, 21, 20], [0, 16, 17, 1, 19, 18],
			[2, 22, 26, 3, 29, 25], [2, 23, 27, 3, 28, 24], [4, 6, 8, 5, 13, 11],
			[4, 7, 9, 5, 12, 10], [6, 16, 25, 13, 19, 26], [7, 17, 24, 12, 18, 27],
			[8, 14, 23, 11, 21, 28], [9, 15, 22, 10, 20, 29],
			[0, 14, 23, 27, 18], [0, 20, 29, 25, 16], [1, 17, 24, 28, 21],
			[1, 19, 26, 22, 15], [2, 22, 10, 12, 24], [2, 25, 13, 11, 23],
			[3, 27, 7, 9, 29], [3, 28, 8, 6, 26], [4, 6, 16, 17, 7],
			[4, 11, 21, 20, 10], [5, 12, 18, 19, 13], [5, 9, 15, 14, 8]]
	},
	Polyhedron{
		name:      'GreatDodecacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.618034
			z: -0.3819660
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: -0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: -0.5801787
			y: 0.0
			z: -0.2216086
		}, Vertex{
			x: -0.5801787
			y: 0.0
			z: 0.2216086
		}, Vertex{
			x: 0.5801787
			y: 0.0
			z: -0.2216086
		}, Vertex{
			x: 0.5801787
			y: 0.0
			z: 0.2216086
		}, Vertex{
			x: 0.0
			y: -0.2216086
			z: -0.5801787
		}, Vertex{
			x: 0.0
			y: -0.2216086
			z: 0.5801787
		}, Vertex{
			x: 0.0
			y: 0.2216086
			z: -0.5801787
		}, Vertex{
			x: 0.0
			y: 0.2216086
			z: 0.5801787
		}, Vertex{
			x: -0.2216086
			y: -0.5801787
			z: 0.0
		}, Vertex{
			x: 0.2216086
			y: -0.5801787
			z: 0.0
		}, Vertex{
			x: -0.2216086
			y: 0.5801787
			z: 0.0
		}, Vertex{
			x: 0.2216086
			y: 0.5801787
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.4606553
			z: 0.2847007
		}, Vertex{
			x: 0.0
			y: -0.4606553
			z: -0.2847007
		}, Vertex{
			x: 0.0
			y: 0.4606553
			z: 0.2847007
		}, Vertex{
			x: 0.0
			y: 0.4606553
			z: -0.2847007
		}, Vertex{
			x: -0.4606553
			y: 0.2847007
			z: 0.0
		}, Vertex{
			x: 0.4606553
			y: 0.2847007
			z: 0.0
		}, Vertex{
			x: -0.4606553
			y: -0.2847007
			z: 0.0
		}, Vertex{
			x: 0.4606553
			y: -0.2847007
			z: 0.0
		}, Vertex{
			x: 0.2847007
			y: 0.0
			z: -0.4606553
		}, Vertex{
			x: 0.2847007
			y: 0.0
			z: 0.4606553
		}, Vertex{
			x: -0.2847007
			y: 0.0
			z: -0.4606553
		}, Vertex{
			x: -0.2847007
			y: 0.0
			z: 0.4606553
		}, Vertex{
			x: 0.3585702
			y: 0.3585702
			z: 0.3585702
		}, Vertex{
			x: 0.3585702
			y: 0.3585702
			z: -0.3585702
		}, Vertex{
			x: -0.3585702
			y: 0.3585702
			z: 0.3585702
		}, Vertex{
			x: -0.3585702
			y: 0.3585702
			z: -0.3585702
		}, Vertex{
			x: 0.3585702
			y: -0.3585702
			z: 0.3585702
		}, Vertex{
			x: 0.3585702
			y: -0.3585702
			z: -0.3585702
		}, Vertex{
			x: -0.3585702
			y: -0.3585702
			z: 0.3585702
		}, Vertex{
			x: -0.3585702
			y: -0.3585702
			z: -0.3585702
		}]
		faces:     [[24, 2, 14, 10], [24, 10, 38, 5], [24, 5, 16, 4],
			[24, 4, 36, 8], [24, 8, 12, 2], [25, 3, 13, 9], [25, 9, 37, 4],
			[25, 4, 17, 5], [25, 5, 39, 11], [25, 11, 15, 3],
			[26, 0, 12, 8], [26, 8, 40, 6], [26, 6, 18, 7], [26, 7, 42, 10],
			[26, 10, 14, 0], [27, 1, 15, 11], [27, 11, 43, 7],
			[27, 7, 19, 6], [27, 6, 41, 9], [27, 9, 13, 1], [28, 0, 16, 5],
			[28, 5, 17, 1], [28, 1, 37, 9], [28, 9, 20, 8], [28, 8, 36, 0],
			[29, 0, 38, 10], [29, 10, 21, 11], [29, 11, 39, 1],
			[29, 1, 17, 4], [29, 4, 16, 0], [30, 2, 40, 8], [30, 8, 22, 9],
			[30, 9, 41, 3], [30, 3, 19, 7], [30, 7, 18, 2], [31, 2, 18, 6],
			[31, 6, 19, 3], [31, 3, 43, 11], [31, 11, 23, 10],
			[31, 10, 42, 2], [32, 0, 36, 4], [32, 4, 20, 9], [32, 9, 22, 6],
			[32, 6, 40, 2], [32, 2, 12, 0], [33, 1, 13, 3], [33, 3, 41, 6],
			[33, 6, 22, 8], [33, 8, 20, 4], [33, 4, 37, 1], [34, 0, 14, 2],
			[34, 2, 42, 7], [34, 7, 23, 11], [34, 11, 21, 5],
			[34, 5, 38, 0], [35, 1, 39, 5], [35, 5, 21, 10], [35, 10, 23, 7],
			[35, 7, 43, 3], [35, 3, 15, 1]]
	},
	Polyhedron{
		name:      'TruncatedOctahedron'
		vertexes_: [Vertex{
			x: 0.7071068
			y: 0.0
			z: 1.414214
		}, Vertex{
			x: 0.7071068
			y: 0.0
			z: -1.414214
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: 1.414214
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: 1.414214
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: -1.414214
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: -1.414214
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.414214
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: 1.414214
			z: -0.7071068
		}, Vertex{
			x: 0.0
			y: -1.414214
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: -1.414214
			z: -0.7071068
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: 1.414214
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: -1.414214
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: 1.414214
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: 1.414214
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: -1.414214
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: -1.414214
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: 0.7071068
			y: 1.414214
			z: 0.0
		}, Vertex{
			x: 0.7071068
			y: -1.414214
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: 1.414214
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: -1.414214
			z: 0.0
		}]
		faces:     [[0, 14, 10, 21, 5, 16], [1, 13, 9, 20, 4, 17],
			[2, 12, 8, 22, 6, 18], [3, 15, 11, 23, 7, 19], [4, 20, 8, 12, 0, 16],
			[5, 21, 11, 15, 1, 17], [7, 23, 10, 14, 2, 18], [6, 22, 9, 13, 3, 19],
			[0, 12, 2, 14], [1, 15, 3, 13], [4, 16, 5, 17], [6, 19, 7, 18],
			[8, 20, 9, 22], [10, 23, 11, 21]]
	},
	Polyhedron{
		name:      'Cuboctahedron'
		vertexes_: [Vertex{
			x: 0.7071068
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: 0.7071068
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: -0.7071068
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: -0.7071068
		}]
		faces:     [[0, 5, 1, 4], [0, 8, 2, 10], [7, 2, 6, 3],
			[7, 11, 5, 10], [9, 1, 11, 3], [9, 6, 8, 4], [0, 4, 8],
			[1, 5, 11], [2, 7, 10], [3, 6, 9], [4, 1, 9], [5, 0, 10],
			[6, 2, 8], [7, 3, 11]]
	},
	Polyhedron{
		name:      'SmallStellatedDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: 0.0
			z: -0.5
		}]
		faces:     [[0, 2, 7, 11, 5], [0, 5, 1, 9, 8], [0, 8, 6, 7, 10],
			[1, 3, 6, 8, 4], [1, 4, 0, 10, 11], [1, 11, 7, 6, 9],
			[2, 0, 4, 9, 6], [2, 6, 3, 11, 10], [2, 10, 5, 4, 8],
			[3, 1, 5, 10, 7], [3, 7, 2, 8, 9], [3, 9, 4, 5, 11]]
	},
	Polyhedron{
		name:      'SmallRetrosnubIcosicosidodecahedron'
		vertexes_: [Vertex{
			x: -0.5768607
			y: 0.0
			z: 0.0666198
		}, Vertex{
			x: -0.5768607
			y: 0.0
			z: -0.0666198
		}, Vertex{
			x: 0.5768607
			y: 0.0
			z: 0.0666198
		}, Vertex{
			x: 0.5768607
			y: 0.0
			z: -0.0666198
		}, Vertex{
			x: 0.0666198
			y: -0.5768607
			z: 0.0
		}, Vertex{
			x: 0.0666198
			y: 0.5768607
			z: 0.0
		}, Vertex{
			x: -0.0666198
			y: -0.5768607
			z: 0.0
		}, Vertex{
			x: -0.0666198
			y: 0.5768607
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.0666198
			z: -0.5768607
		}, Vertex{
			x: 0.0
			y: 0.0666198
			z: 0.5768607
		}, Vertex{
			x: 0.0
			y: -0.0666198
			z: -0.5768607
		}, Vertex{
			x: 0.0
			y: -0.0666198
			z: 0.5768607
		}, Vertex{
			x: -0.2678437
			y: 0.5
			z: -0.1243632
		}, Vertex{
			x: -0.2678437
			y: 0.5
			z: 0.1243632
		}, Vertex{
			x: -0.2678437
			y: -0.5
			z: -0.1243632
		}, Vertex{
			x: -0.2678437
			y: -0.5
			z: 0.1243632
		}, Vertex{
			x: 0.2678437
			y: 0.5
			z: -0.1243632
		}, Vertex{
			x: 0.2678437
			y: 0.5
			z: 0.1243632
		}, Vertex{
			x: 0.2678437
			y: -0.5
			z: -0.1243632
		}, Vertex{
			x: 0.2678437
			y: -0.5
			z: 0.1243632
		}, Vertex{
			x: -0.1243632
			y: -0.2678437
			z: 0.5
		}, Vertex{
			x: -0.1243632
			y: -0.2678437
			z: -0.5
		}, Vertex{
			x: -0.1243632
			y: 0.2678437
			z: 0.5
		}, Vertex{
			x: -0.1243632
			y: 0.2678437
			z: -0.5
		}, Vertex{
			x: 0.1243632
			y: -0.2678437
			z: 0.5
		}, Vertex{
			x: 0.1243632
			y: -0.2678437
			z: -0.5
		}, Vertex{
			x: 0.1243632
			y: 0.2678437
			z: 0.5
		}, Vertex{
			x: 0.1243632
			y: 0.2678437
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.1243632
			z: -0.2678437
		}, Vertex{
			x: 0.5
			y: -0.1243632
			z: 0.2678437
		}, Vertex{
			x: 0.5
			y: 0.1243632
			z: -0.2678437
		}, Vertex{
			x: 0.5
			y: 0.1243632
			z: 0.2678437
		}, Vertex{
			x: -0.5
			y: -0.1243632
			z: -0.2678437
		}, Vertex{
			x: -0.5
			y: -0.1243632
			z: 0.2678437
		}, Vertex{
			x: -0.5
			y: 0.1243632
			z: -0.2678437
		}, Vertex{
			x: -0.5
			y: 0.1243632
			z: 0.2678437
		}, Vertex{
			x: 0.309017
			y: -0.4333802
			z: 0.2321563
		}, Vertex{
			x: 0.309017
			y: -0.4333802
			z: -0.2321563
		}, Vertex{
			x: 0.309017
			y: 0.4333802
			z: 0.2321563
		}, Vertex{
			x: 0.309017
			y: 0.4333802
			z: -0.2321563
		}, Vertex{
			x: -0.309017
			y: -0.4333802
			z: 0.2321563
		}, Vertex{
			x: -0.309017
			y: -0.4333802
			z: -0.2321563
		}, Vertex{
			x: -0.309017
			y: 0.4333802
			z: 0.2321563
		}, Vertex{
			x: -0.309017
			y: 0.4333802
			z: -0.2321563
		}, Vertex{
			x: 0.2321563
			y: 0.309017
			z: -0.4333802
		}, Vertex{
			x: 0.2321563
			y: 0.309017
			z: 0.4333802
		}, Vertex{
			x: 0.2321563
			y: -0.309017
			z: -0.4333802
		}, Vertex{
			x: 0.2321563
			y: -0.309017
			z: 0.4333802
		}, Vertex{
			x: -0.2321563
			y: 0.309017
			z: -0.4333802
		}, Vertex{
			x: -0.2321563
			y: 0.309017
			z: 0.4333802
		}, Vertex{
			x: -0.2321563
			y: -0.309017
			z: -0.4333802
		}, Vertex{
			x: -0.2321563
			y: -0.309017
			z: 0.4333802
		}, Vertex{
			x: -0.4333802
			y: 0.2321563
			z: 0.309017
		}, Vertex{
			x: -0.4333802
			y: 0.2321563
			z: -0.309017
		}, Vertex{
			x: -0.4333802
			y: -0.2321563
			z: 0.309017
		}, Vertex{
			x: -0.4333802
			y: -0.2321563
			z: -0.309017
		}, Vertex{
			x: 0.4333802
			y: 0.2321563
			z: 0.309017
		}, Vertex{
			x: 0.4333802
			y: 0.2321563
			z: -0.309017
		}, Vertex{
			x: 0.4333802
			y: -0.2321563
			z: 0.309017
		}, Vertex{
			x: 0.4333802
			y: -0.2321563
			z: -0.309017
		}]
		faces:     [[0, 46, 12, 14, 44], [1, 45, 15, 13, 47],
			[2, 48, 18, 16, 50], [3, 51, 17, 19, 49], [4, 53, 20, 21, 52],
			[5, 54, 23, 22, 55], [6, 56, 25, 24, 57], [7, 59, 26, 27, 58],
			[8, 40, 28, 32, 36], [9, 37, 33, 29, 41], [10, 38, 34, 30, 42],
			[11, 43, 31, 35, 39], [0, 16, 18], [1, 19, 17], [2, 14, 12],
			[3, 13, 15], [4, 22, 23], [5, 21, 20], [6, 27, 26],
			[7, 24, 25], [8, 29, 33], [9, 32, 28], [10, 35, 31],
			[11, 30, 34], [12, 28, 40], [13, 41, 29], [14, 42, 30],
			[15, 31, 43], [16, 36, 32], [17, 33, 37], [18, 34, 38],
			[19, 39, 35], [20, 12, 46], [21, 47, 13], [22, 44, 14],
			[23, 15, 45], [24, 50, 16], [25, 17, 51], [26, 18, 48],
			[27, 49, 19], [28, 20, 53], [29, 52, 21], [30, 55, 22],
			[31, 23, 54], [32, 57, 24], [33, 25, 56], [34, 26, 59],
			[35, 58, 27], [36, 0, 44], [37, 45, 1], [38, 46, 0],
			[39, 1, 47], [40, 48, 2], [41, 3, 49], [42, 2, 50],
			[43, 51, 3], [44, 4, 52], [45, 53, 4], [46, 54, 5],
			[47, 5, 55], [48, 56, 6], [49, 6, 57], [50, 7, 58],
			[51, 59, 7], [52, 8, 36], [53, 37, 9], [54, 38, 10],
			[55, 11, 39], [56, 40, 8], [57, 9, 41], [58, 10, 42],
			[59, 43, 11], [0, 18, 38], [0, 36, 16], [1, 17, 37],
			[1, 39, 19], [2, 12, 40], [2, 42, 14], [3, 15, 43],
			[3, 41, 13], [21, 5, 47], [21, 13, 29], [22, 4, 44],
			[22, 14, 30], [25, 33, 17], [25, 51, 7], [26, 34, 18],
			[26, 48, 6], [28, 12, 20], [28, 53, 9], [31, 15, 23],
			[31, 54, 10], [32, 9, 57], [32, 24, 16], [35, 10, 58],
			[35, 27, 19], [45, 4, 23], [45, 37, 53], [46, 5, 20],
			[46, 38, 54], [49, 27, 6], [49, 57, 41], [50, 24, 7],
			[50, 58, 42], [52, 29, 8], [52, 36, 44], [55, 30, 11],
			[55, 39, 47], [56, 8, 33], [56, 48, 40], [59, 11, 34],
			[59, 51, 43]]
	},
	Polyhedron{
		name:      'SmallRhombihexahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: -0.5
		}]
		faces:     [[0, 2, 18, 19, 3, 1, 17, 16], [0, 8, 9, 1, 5, 13, 12, 4],
			[14, 15, 7, 3, 11, 10, 2, 6], [14, 22, 18, 10, 8, 16, 20, 12],
			[21, 5, 7, 23, 22, 6, 4, 20], [21, 17, 9, 11, 19, 23, 15, 13],
			[0, 2, 10, 8], [0, 16, 20, 4], [7, 3, 19, 23], [7, 15, 13, 5],
			[11, 3, 1, 9], [11, 10, 18, 19], [12, 14, 6, 4], [12, 20, 21, 13],
			[17, 1, 5, 21], [17, 16, 8, 9], [22, 14, 15, 23],
			[22, 18, 2, 6]]
	},
	Polyhedron{
		name:      'GreatIcosihemidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: -0.309017
			z: 0.5
		}]
		faces:     [[0, 6, 22, 23, 7, 1, 13, 29, 28, 12], [0, 8, 24, 25, 9, 1, 11, 27, 26, 10],
			[2, 14, 6, 10, 18, 3, 21, 13, 9, 17], [2, 15, 7, 11, 19, 3, 20, 12, 8, 16],
			[4, 22, 14, 16, 24, 5, 29, 21, 19, 27], [4, 23, 15, 17, 25, 5, 28, 20, 18, 26],
			[0, 6, 10], [0, 12, 8], [1, 9, 13], [1, 11, 7], [14, 16, 2],
			[14, 22, 6], [17, 15, 2], [17, 25, 9], [19, 21, 3],
			[19, 27, 11], [20, 18, 3], [20, 28, 12], [23, 4, 22],
			[23, 15, 7], [24, 5, 25], [24, 16, 8], [26, 4, 27],
			[26, 18, 10], [29, 5, 28], [29, 21, 13]]
	},
	Polyhedron{
		name:      'Octahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: 0.0
		}]
		faces:     [[0, 2, 4], [0, 4, 3], [0, 3, 5], [0, 5, 2],
			[1, 2, 5], [1, 5, 3], [1, 3, 4], [1, 4, 2]]
	},
	Polyhedron{
		name:      'GreatStellatedDodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: 0.0
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: 0.0
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: 0.0
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: 0.0
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: 0.0
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: -0.309017
			z: -0.309017
		}, Vertex{
			x: -0.309017
			y: -0.309017
			z: 0.309017
		}, Vertex{
			x: 0.309017
			y: -0.309017
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: -0.309017
			z: 0.309017
		}, Vertex{
			x: -0.309017
			y: 0.309017
			z: -0.309017
		}, Vertex{
			x: -0.309017
			y: 0.309017
			z: 0.309017
		}, Vertex{
			x: 0.309017
			y: 0.309017
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: 0.309017
			z: 0.309017
		}]
		faces:     [[0, 2, 14, 4, 12], [0, 12, 8, 10, 16], [0, 16, 6, 18, 2],
			[7, 6, 16, 10, 17], [7, 17, 1, 3, 19], [7, 19, 11, 18, 6],
			[9, 11, 19, 3, 15], [9, 15, 5, 4, 14], [9, 14, 2, 18, 11],
			[13, 1, 17, 10, 8], [13, 8, 12, 4, 5], [13, 5, 15, 3, 1]]
	},
	Polyhedron{
		name:      'Rhombidodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.1909830
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: 1.0
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: -1.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: 1.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: -1.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: 1.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: -1.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: 1.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: 1.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: 1.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: 1.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: -1.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: -1.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: -1.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: -1.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: 1.0
			z: -0.309017
		}, Vertex{
			x: 0.809017
			y: -1.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: -1.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: 1.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: 1.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: -1.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: -1.0
			z: -0.309017
		}]
		faces:     [[0, 40, 24, 26, 42], [1, 43, 27, 25, 41],
			[2, 38, 22, 20, 36], [3, 37, 21, 23, 39], [4, 46, 30, 31, 47],
			[5, 45, 29, 28, 44], [6, 51, 35, 34, 50], [7, 48, 32, 33, 49],
			[8, 53, 13, 17, 57], [9, 56, 16, 12, 52], [10, 59, 19, 15, 55],
			[11, 54, 14, 18, 58], [0, 46, 12, 14, 44], [1, 45, 15, 13, 47],
			[2, 48, 18, 16, 50], [3, 51, 17, 19, 49], [4, 53, 20, 21, 52],
			[5, 54, 23, 22, 55], [6, 56, 25, 24, 57], [7, 59, 26, 27, 58],
			[8, 40, 28, 32, 36], [9, 37, 33, 29, 41], [10, 38, 34, 30, 42],
			[11, 43, 31, 35, 39], [0, 42, 30, 46], [0, 44, 28, 40],
			[1, 41, 29, 45], [1, 47, 31, 43], [3, 39, 35, 51],
			[3, 49, 33, 37], [5, 44, 14, 54], [5, 55, 15, 45],
			[6, 50, 16, 56], [6, 57, 17, 51], [7, 49, 19, 59],
			[7, 58, 18, 48], [8, 36, 20, 53], [8, 57, 24, 40],
			[9, 41, 25, 56], [9, 52, 21, 37], [11, 39, 23, 54],
			[11, 58, 27, 43], [12, 16, 18, 14], [12, 46, 4, 52],
			[13, 15, 19, 17], [13, 53, 4, 47], [22, 23, 21, 20],
			[22, 38, 10, 55], [26, 24, 25, 27], [26, 59, 10, 42],
			[32, 28, 29, 33], [32, 48, 2, 36], [34, 35, 31, 30],
			[34, 38, 2, 50]]
	},
	Polyhedron{
		name:      'Icosidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: -1.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: 1.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: -1.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: 1.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: 1.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: 1.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: -1.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: -1.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: -1.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: 1.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: 1.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: -1.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: -1.309017
			z: -0.5
		}]
		faces:     [[0, 8, 16, 14, 6], [0, 10, 18, 20, 12], [1, 7, 15, 17, 9],
			[1, 13, 21, 19, 11], [2, 15, 23, 22, 14], [2, 16, 24, 25, 17],
			[3, 18, 26, 27, 19], [3, 21, 29, 28, 20], [4, 23, 7, 11, 27],
			[4, 26, 10, 6, 22], [5, 24, 8, 12, 28], [5, 29, 13, 9, 25],
			[0, 6, 10], [0, 12, 8], [1, 9, 13], [1, 11, 7], [2, 14, 16],
			[2, 17, 15], [3, 19, 21], [3, 20, 18], [4, 22, 23],
			[4, 27, 26], [5, 25, 24], [5, 28, 29], [6, 14, 22],
			[7, 23, 15], [8, 24, 16], [9, 17, 25], [10, 26, 18],
			[11, 19, 27], [12, 20, 28], [13, 29, 21]]
	},
	Polyhedron{
		name:      'SmallStellapentakisDodecahedron'
		vertexes_: [Vertex{
			x: 1.809017
			y: 0.0
			z: 2.927051
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -2.927051
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 2.927051
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -2.927051
		}, Vertex{
			x: 2.927051
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 2.927051
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -2.927051
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -2.927051
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.927051
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 2.927051
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -2.927051
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -2.927051
			z: -1.809017
		}, Vertex{
			x: 0.9549151
			y: 0.0
			z: 1.545085
		}, Vertex{
			x: 0.9549151
			y: 0.0
			z: -1.545085
		}, Vertex{
			x: -0.9549151
			y: 0.0
			z: 1.545085
		}, Vertex{
			x: -0.9549151
			y: 0.0
			z: -1.545085
		}, Vertex{
			x: 1.545085
			y: 0.9549151
			z: 0.0
		}, Vertex{
			x: 1.545085
			y: -0.9549151
			z: 0.0
		}, Vertex{
			x: -1.545085
			y: 0.9549151
			z: 0.0
		}, Vertex{
			x: -1.545085
			y: -0.9549151
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.545085
			z: 0.9549151
		}, Vertex{
			x: 0.0
			y: 1.545085
			z: -0.9549151
		}, Vertex{
			x: 0.0
			y: -1.545085
			z: 0.9549151
		}, Vertex{
			x: 0.0
			y: -1.545085
			z: -0.9549151
		}]
		faces:     [[12, 2, 5], [12, 5, 8], [12, 8, 10], [12, 10, 4],
			[12, 4, 2], [13, 3, 4], [13, 4, 11], [13, 11, 9],
			[13, 9, 5], [13, 5, 3], [14, 0, 6], [14, 6, 10], [14, 10, 8],
			[14, 8, 7], [14, 7, 0], [15, 1, 7], [15, 7, 9], [15, 9, 11],
			[15, 11, 6], [15, 6, 1], [16, 0, 1], [16, 1, 8], [16, 8, 5],
			[16, 5, 9], [16, 9, 0], [17, 1, 0], [17, 0, 11], [17, 11, 4],
			[17, 4, 10], [17, 10, 1], [18, 3, 2], [18, 2, 9],
			[18, 9, 7], [18, 7, 8], [18, 8, 3], [19, 2, 3], [19, 3, 10],
			[19, 10, 6], [19, 6, 11], [19, 11, 2], [20, 0, 9],
			[20, 9, 2], [20, 2, 4], [20, 4, 6], [20, 6, 0], [21, 1, 6],
			[21, 6, 4], [21, 4, 3], [21, 3, 8], [21, 8, 1], [22, 0, 7],
			[22, 7, 5], [22, 5, 2], [22, 2, 11], [22, 11, 0],
			[23, 1, 10], [23, 10, 3], [23, 3, 5], [23, 5, 7],
			[23, 7, 1]]
	},
	Polyhedron{
		name:      'GreatStellatedTruncatedDodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.0
			z: -0.4270510
		}, Vertex{
			x: 0.5
			y: 0.0
			z: 0.4270510
		}, Vertex{
			x: -0.5
			y: 0.0
			z: -0.4270510
		}, Vertex{
			x: -0.5
			y: 0.0
			z: 0.4270510
		}, Vertex{
			x: 0.0
			y: -0.4270510
			z: 0.5
		}, Vertex{
			x: 0.0
			y: -0.4270510
			z: -0.5
		}, Vertex{
			x: 0.0
			y: 0.4270510
			z: 0.5
		}, Vertex{
			x: 0.0
			y: 0.4270510
			z: -0.5
		}, Vertex{
			x: -0.4270510
			y: 0.5
			z: 0.0
		}, Vertex{
			x: 0.4270510
			y: 0.5
			z: 0.0
		}, Vertex{
			x: -0.4270510
			y: -0.5
			z: 0.0
		}, Vertex{
			x: 0.4270510
			y: -0.5
			z: 0.0
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: 0.3819660
		}, Vertex{
			x: 0.1909830
			y: 0.5
			z: -0.3819660
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: 0.3819660
		}, Vertex{
			x: -0.1909830
			y: 0.5
			z: -0.3819660
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: 0.3819660
		}, Vertex{
			x: 0.1909830
			y: -0.5
			z: -0.3819660
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: 0.3819660
		}, Vertex{
			x: -0.1909830
			y: -0.5
			z: -0.3819660
		}, Vertex{
			x: 0.5
			y: 0.3819660
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: 0.3819660
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: 0.3819660
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: 0.3819660
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: -0.3819660
			z: 0.1909830
		}, Vertex{
			x: 0.5
			y: -0.3819660
			z: -0.1909830
		}, Vertex{
			x: -0.5
			y: -0.3819660
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: -0.3819660
			z: -0.1909830
		}, Vertex{
			x: 0.3819660
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: 0.3819660
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: -0.3819660
			y: 0.1909830
			z: 0.5
		}, Vertex{
			x: -0.3819660
			y: 0.1909830
			z: -0.5
		}, Vertex{
			x: 0.3819660
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: 0.3819660
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: -0.3819660
			y: -0.1909830
			z: 0.5
		}, Vertex{
			x: -0.3819660
			y: -0.1909830
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: 0.1909830
			z: -0.1180340
		}, Vertex{
			x: -0.618034
			y: 0.1909830
			z: 0.1180340
		}, Vertex{
			x: 0.618034
			y: 0.1909830
			z: -0.1180340
		}, Vertex{
			x: 0.618034
			y: 0.1909830
			z: 0.1180340
		}, Vertex{
			x: -0.618034
			y: -0.1909830
			z: -0.1180340
		}, Vertex{
			x: -0.618034
			y: -0.1909830
			z: 0.1180340
		}, Vertex{
			x: 0.618034
			y: -0.1909830
			z: -0.1180340
		}, Vertex{
			x: 0.618034
			y: -0.1909830
			z: 0.1180340
		}, Vertex{
			x: 0.1909830
			y: -0.1180340
			z: -0.618034
		}, Vertex{
			x: 0.1909830
			y: -0.1180340
			z: 0.618034
		}, Vertex{
			x: -0.1909830
			y: -0.1180340
			z: -0.618034
		}, Vertex{
			x: -0.1909830
			y: -0.1180340
			z: 0.618034
		}, Vertex{
			x: 0.1909830
			y: 0.1180340
			z: -0.618034
		}, Vertex{
			x: 0.1909830
			y: 0.1180340
			z: 0.618034
		}, Vertex{
			x: -0.1909830
			y: 0.1180340
			z: -0.618034
		}, Vertex{
			x: -0.1909830
			y: 0.1180340
			z: 0.618034
		}, Vertex{
			x: -0.1180340
			y: -0.618034
			z: 0.1909830
		}, Vertex{
			x: -0.1180340
			y: -0.618034
			z: -0.1909830
		}, Vertex{
			x: 0.1180340
			y: -0.618034
			z: 0.1909830
		}, Vertex{
			x: 0.1180340
			y: -0.618034
			z: -0.1909830
		}, Vertex{
			x: -0.1180340
			y: 0.618034
			z: 0.1909830
		}, Vertex{
			x: -0.1180340
			y: 0.618034
			z: -0.1909830
		}, Vertex{
			x: 0.1180340
			y: 0.618034
			z: 0.1909830
		}, Vertex{
			x: 0.1180340
			y: 0.618034
			z: -0.1909830
		}]
		faces:     [[0, 2, 14, 38, 46, 22, 20, 44, 36, 12], [1, 3, 19, 43, 51, 27, 25, 49, 41, 17],
			[2, 0, 16, 40, 48, 24, 26, 50, 42, 18], [3, 1, 13, 37, 45, 21, 23, 47, 39, 15],
			[4, 5, 21, 45, 53, 29, 28, 52, 44, 20], [5, 4, 22, 46, 54, 30, 31, 55, 47, 23],
			[6, 7, 27, 51, 59, 35, 34, 58, 50, 26], [7, 6, 24, 48, 56, 32, 33, 57, 49, 25],
			[8, 10, 32, 56, 40, 16, 12, 36, 52, 28], [9, 11, 35, 59, 43, 19, 15, 39, 55, 31],
			[10, 8, 29, 53, 37, 13, 17, 41, 57, 33], [11, 9, 30, 54, 38, 14, 18, 42, 58, 34],
			[0, 12, 16], [1, 17, 13], [2, 18, 14], [3, 15, 19],
			[4, 20, 22], [5, 23, 21], [6, 26, 24], [7, 25, 27],
			[8, 28, 29], [9, 31, 30], [10, 33, 32], [11, 34, 35],
			[36, 44, 52], [37, 53, 45], [38, 54, 46], [39, 47, 55],
			[40, 56, 48], [41, 49, 57], [42, 50, 58], [43, 59, 51]]
	},
	Polyhedron{
		name:      'Icosahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.0
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: 0.0
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: 0.0
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: 0.0
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: 0.0
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: 0.0
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: 0.0
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: 0.0
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: 0.0
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: 0.0
			y: -0.809017
			z: -0.5
		}]
		faces:     [[0, 2, 10], [0, 10, 5], [0, 5, 4], [0, 4, 8],
			[0, 8, 2], [3, 1, 11], [3, 11, 7], [3, 7, 6], [3, 6, 9],
			[3, 9, 1], [2, 6, 7], [2, 7, 10], [10, 7, 11], [10, 11, 5],
			[5, 11, 1], [5, 1, 4], [4, 1, 9], [4, 9, 8], [8, 9, 6],
			[8, 6, 2]]
	},
	Polyhedron{
		name:      'PentagonalHexecontahedron(laevo}'
		vertexes_: [Vertex{
			x: -0.1928937
			y: -0.2184834
			z: -2.097054
		}, Vertex{
			x: -0.1928937
			y: 0.2184834
			z: 2.097054
		}, Vertex{
			x: 0.1928937
			y: 0.2184834
			z: -2.097054
		}, Vertex{
			x: 0.1928937
			y: -0.2184834
			z: 2.097054
		}, Vertex{
			x: -2.097054
			y: -0.1928937
			z: -0.2184834
		}, Vertex{
			x: -2.097054
			y: 0.1928937
			z: 0.2184834
		}, Vertex{
			x: 2.097054
			y: 0.1928937
			z: -0.2184834
		}, Vertex{
			x: 2.097054
			y: -0.1928937
			z: 0.2184834
		}, Vertex{
			x: -0.2184834
			y: -2.097054
			z: -0.1928937
		}, Vertex{
			x: -0.2184834
			y: 2.097054
			z: 0.1928937
		}, Vertex{
			x: 0.2184834
			y: 2.097054
			z: -0.1928937
		}, Vertex{
			x: 0.2184834
			y: -2.097054
			z: 0.1928937
		}, Vertex{
			x: 0.0
			y: -0.7554672
			z: -1.977839
		}, Vertex{
			x: 0.0
			y: -0.7554672
			z: 1.977839
		}, Vertex{
			x: 0.0
			y: 0.7554672
			z: -1.977839
		}, Vertex{
			x: 0.0
			y: 0.7554672
			z: 1.977839
		}, Vertex{
			x: -1.977839
			y: 0.0
			z: -0.7554672
		}, Vertex{
			x: -1.977839
			y: 0.0
			z: 0.7554672
		}, Vertex{
			x: 1.977839
			y: 0.0
			z: -0.7554672
		}, Vertex{
			x: 1.977839
			y: 0.0
			z: 0.7554672
		}, Vertex{
			x: -0.7554672
			y: -1.977839
			z: 0.0
		}, Vertex{
			x: -0.7554672
			y: 1.977839
			z: 0.0
		}, Vertex{
			x: 0.7554672
			y: -1.977839
			z: 0.0
		}, Vertex{
			x: 0.7554672
			y: 1.977839
			z: 0.0
		}, Vertex{
			x: -1.167123
			y: 0.0
			z: -1.888445
		}, Vertex{
			x: -1.167123
			y: 0.0
			z: 1.888445
		}, Vertex{
			x: 1.167123
			y: 0.0
			z: -1.888445
		}, Vertex{
			x: 1.167123
			y: 0.0
			z: 1.888445
		}, Vertex{
			x: -1.888445
			y: -1.167123
			z: 0.0
		}, Vertex{
			x: -1.888445
			y: 1.167123
			z: 0.0
		}, Vertex{
			x: 1.888445
			y: -1.167123
			z: 0.0
		}, Vertex{
			x: 1.888445
			y: 1.167123
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.888445
			z: -1.167123
		}, Vertex{
			x: 0.0
			y: -1.888445
			z: 1.167123
		}, Vertex{
			x: 0.0
			y: 1.888445
			z: -1.167123
		}, Vertex{
			x: 0.0
			y: 1.888445
			z: 1.167123
		}, Vertex{
			x: -0.5677154
			y: 0.8249576
			z: -1.865401
		}, Vertex{
			x: -0.5677154
			y: -0.8249576
			z: 1.865401
		}, Vertex{
			x: 0.5677154
			y: -0.8249576
			z: -1.865401
		}, Vertex{
			x: 0.5677154
			y: 0.8249576
			z: 1.865401
		}, Vertex{
			x: -1.865401
			y: 0.5677154
			z: -0.8249576
		}, Vertex{
			x: -1.865401
			y: -0.5677154
			z: 0.8249576
		}, Vertex{
			x: 1.865401
			y: -0.5677154
			z: -0.8249576
		}, Vertex{
			x: 1.865401
			y: 0.5677154
			z: 0.8249576
		}, Vertex{
			x: -0.8249576
			y: 1.865401
			z: -0.5677154
		}, Vertex{
			x: -0.8249576
			y: -1.865401
			z: 0.5677154
		}, Vertex{
			x: 0.8249576
			y: -1.865401
			z: -0.5677154
		}, Vertex{
			x: 0.8249576
			y: 1.865401
			z: 0.5677154
		}, Vertex{
			x: -0.3748217
			y: -1.137066
			z: -1.746187
		}, Vertex{
			x: -0.3748217
			y: 1.137066
			z: 1.746187
		}, Vertex{
			x: 0.3748217
			y: 1.137066
			z: -1.746187
		}, Vertex{
			x: 0.3748217
			y: -1.137066
			z: 1.746187
		}, Vertex{
			x: -1.746187
			y: -0.3748217
			z: -1.137066
		}, Vertex{
			x: -1.746187
			y: 0.3748217
			z: 1.137066
		}, Vertex{
			x: 1.746187
			y: 0.3748217
			z: -1.137066
		}, Vertex{
			x: 1.746187
			y: -0.3748217
			z: 1.137066
		}, Vertex{
			x: -1.137066
			y: -1.746187
			z: -0.3748217
		}, Vertex{
			x: -1.137066
			y: 1.746187
			z: 0.3748217
		}, Vertex{
			x: 1.137066
			y: 1.746187
			z: -0.3748217
		}, Vertex{
			x: 1.137066
			y: -1.746187
			z: 0.3748217
		}, Vertex{
			x: -0.9212289
			y: -0.9599877
			z: -1.646918
		}, Vertex{
			x: -0.9212289
			y: 0.9599877
			z: 1.646918
		}, Vertex{
			x: 0.9212289
			y: 0.9599877
			z: -1.646918
		}, Vertex{
			x: 0.9212289
			y: -0.9599877
			z: 1.646918
		}, Vertex{
			x: -1.646918
			y: -0.9212289
			z: -0.9599877
		}, Vertex{
			x: -1.646918
			y: 0.9212289
			z: 0.9599877
		}, Vertex{
			x: 1.646918
			y: 0.9212289
			z: -0.9599877
		}, Vertex{
			x: 1.646918
			y: -0.9212289
			z: 0.9599877
		}, Vertex{
			x: -0.9599877
			y: -1.646918
			z: -0.9212289
		}, Vertex{
			x: -0.9599877
			y: 1.646918
			z: 0.9212289
		}, Vertex{
			x: 0.9599877
			y: 1.646918
			z: -0.9212289
		}, Vertex{
			x: 0.9599877
			y: -1.646918
			z: 0.9212289
		}, Vertex{
			x: -0.7283352
			y: 1.272096
			z: -1.527703
		}, Vertex{
			x: -0.7283352
			y: -1.272096
			z: 1.527703
		}, Vertex{
			x: 0.7283352
			y: -1.272096
			z: -1.527703
		}, Vertex{
			x: 0.7283352
			y: 1.272096
			z: 1.527703
		}, Vertex{
			x: -1.527703
			y: 0.7283352
			z: -1.272096
		}, Vertex{
			x: -1.527703
			y: -0.7283352
			z: 1.272096
		}, Vertex{
			x: 1.527703
			y: -0.7283352
			z: -1.272096
		}, Vertex{
			x: 1.527703
			y: 0.7283352
			z: 1.272096
		}, Vertex{
			x: -1.272096
			y: 1.527703
			z: -0.7283352
		}, Vertex{
			x: -1.272096
			y: -1.527703
			z: 0.7283352
		}, Vertex{
			x: 1.272096
			y: -1.527703
			z: -0.7283352
		}, Vertex{
			x: 1.272096
			y: 1.527703
			z: 0.7283352
		}, Vertex{
			x: -1.222372
			y: -1.222372
			z: -1.222372
		}, Vertex{
			x: -1.222372
			y: -1.222372
			z: 1.222372
		}, Vertex{
			x: -1.222372
			y: 1.222372
			z: -1.222372
		}, Vertex{
			x: -1.222372
			y: 1.222372
			z: 1.222372
		}, Vertex{
			x: 1.222372
			y: -1.222372
			z: -1.222372
		}, Vertex{
			x: 1.222372
			y: -1.222372
			z: 1.222372
		}, Vertex{
			x: 1.222372
			y: 1.222372
			z: -1.222372
		}, Vertex{
			x: 1.222372
			y: 1.222372
			z: 1.222372
		}]
		faces:     [[24, 36, 14, 2, 0], [24, 76, 86, 72, 36],
			[24, 52, 16, 40, 76], [24, 60, 84, 64, 52], [24, 0, 12, 48, 60],
			[25, 37, 13, 3, 1], [25, 77, 85, 73, 37], [25, 53, 17, 41, 77],
			[25, 61, 87, 65, 53], [25, 1, 15, 49, 61], [26, 38, 12, 0, 2],
			[26, 78, 88, 74, 38], [26, 54, 18, 42, 78], [26, 62, 90, 66, 54],
			[26, 2, 14, 50, 62], [27, 39, 15, 1, 3], [27, 79, 91, 75, 39],
			[27, 55, 19, 43, 79], [27, 63, 89, 67, 55], [27, 3, 13, 51, 63],
			[28, 41, 17, 5, 4], [28, 81, 85, 77, 41], [28, 56, 20, 45, 81],
			[28, 64, 84, 68, 56], [28, 4, 16, 52, 64], [29, 40, 16, 4, 5],
			[29, 80, 86, 76, 40], [29, 57, 21, 44, 80], [29, 65, 87, 69, 57],
			[29, 5, 17, 53, 65], [30, 42, 18, 6, 7], [30, 82, 88, 78, 42],
			[30, 59, 22, 46, 82], [30, 67, 89, 71, 59], [30, 7, 19, 55, 67],
			[31, 43, 19, 7, 6], [31, 83, 91, 79, 43], [31, 58, 23, 47, 83],
			[31, 66, 90, 70, 58], [31, 6, 18, 54, 66], [32, 46, 22, 11, 8],
			[32, 74, 88, 82, 46], [32, 48, 12, 38, 74], [32, 68, 84, 60, 48],
			[32, 8, 20, 56, 68], [33, 45, 20, 8, 11], [33, 73, 85, 81, 45],
			[33, 51, 13, 37, 73], [33, 71, 89, 63, 51], [33, 11, 22, 59, 71],
			[34, 44, 21, 9, 10], [34, 72, 86, 80, 44], [34, 50, 14, 36, 72],
			[34, 70, 90, 62, 50], [34, 10, 23, 58, 70], [35, 47, 23, 10, 9],
			[35, 75, 91, 83, 47], [35, 49, 15, 39, 75], [35, 69, 87, 61, 49],
			[35, 9, 21, 57, 69]]
	},
	Polyhedron{
		name:      'TetradyakisHexahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 7.242641
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -7.242641
		}, Vertex{
			x: 7.242641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -7.242641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 7.242641
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -7.242641
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.242641
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.242641
		}, Vertex{
			x: 1.242641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.242641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.242641
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.242641
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: 1.0
			y: -1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: 1.0
			z: -1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: 1.0
		}, Vertex{
			x: -1.0
			y: -1.0
			z: -1.0
		}]
		faces:     [[0, 8, 13], [0, 13, 10], [0, 10, 17], [0, 17, 9],
			[0, 9, 19], [0, 19, 11], [0, 11, 15], [0, 15, 8],
			[1, 8, 14], [1, 14, 11], [1, 11, 18], [1, 18, 9],
			[1, 9, 16], [1, 16, 10], [1, 10, 12], [1, 12, 8],
			[2, 6, 18], [2, 18, 11], [2, 11, 19], [2, 19, 7],
			[2, 7, 17], [2, 17, 10], [2, 10, 16], [2, 16, 6],
			[3, 6, 12], [3, 12, 10], [3, 10, 13], [3, 13, 7],
			[3, 7, 15], [3, 15, 11], [3, 11, 14], [3, 14, 6],
			[4, 6, 14], [4, 14, 8], [4, 8, 15], [4, 15, 7], [4, 7, 19],
			[4, 19, 9], [4, 9, 18], [4, 18, 6], [5, 6, 16], [5, 16, 9],
			[5, 9, 17], [5, 17, 7], [5, 7, 13], [5, 13, 8], [5, 8, 12],
			[5, 12, 6]]
	},
	Polyhedron{
		name:      'TruncatedIcosahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.0
			z: 2.427051
		}, Vertex{
			x: 0.5
			y: 0.0
			z: -2.427051
		}, Vertex{
			x: -0.5
			y: 0.0
			z: 2.427051
		}, Vertex{
			x: -0.5
			y: 0.0
			z: -2.427051
		}, Vertex{
			x: 2.427051
			y: 0.5
			z: 0.0
		}, Vertex{
			x: 2.427051
			y: -0.5
			z: 0.0
		}, Vertex{
			x: -2.427051
			y: 0.5
			z: 0.0
		}, Vertex{
			x: -2.427051
			y: -0.5
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.427051
			z: 0.5
		}, Vertex{
			x: 0.0
			y: 2.427051
			z: -0.5
		}, Vertex{
			x: 0.0
			y: -2.427051
			z: 0.5
		}, Vertex{
			x: 0.0
			y: -2.427051
			z: -0.5
		}, Vertex{
			x: 1.0
			y: 0.809017
			z: 2.118034
		}, Vertex{
			x: 1.0
			y: 0.809017
			z: -2.118034
		}, Vertex{
			x: 1.0
			y: -0.809017
			z: 2.118034
		}, Vertex{
			x: 1.0
			y: -0.809017
			z: -2.118034
		}, Vertex{
			x: -1.0
			y: 0.809017
			z: 2.118034
		}, Vertex{
			x: -1.0
			y: 0.809017
			z: -2.118034
		}, Vertex{
			x: -1.0
			y: -0.809017
			z: 2.118034
		}, Vertex{
			x: -1.0
			y: -0.809017
			z: -2.118034
		}, Vertex{
			x: 2.118034
			y: 1.0
			z: 0.809017
		}, Vertex{
			x: 2.118034
			y: 1.0
			z: -0.809017
		}, Vertex{
			x: 2.118034
			y: -1.0
			z: 0.809017
		}, Vertex{
			x: 2.118034
			y: -1.0
			z: -0.809017
		}, Vertex{
			x: -2.118034
			y: 1.0
			z: 0.809017
		}, Vertex{
			x: -2.118034
			y: 1.0
			z: -0.809017
		}, Vertex{
			x: -2.118034
			y: -1.0
			z: 0.809017
		}, Vertex{
			x: -2.118034
			y: -1.0
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 2.118034
			z: 1.0
		}, Vertex{
			x: 0.809017
			y: 2.118034
			z: -1.0
		}, Vertex{
			x: 0.809017
			y: -2.118034
			z: 1.0
		}, Vertex{
			x: 0.809017
			y: -2.118034
			z: -1.0
		}, Vertex{
			x: -0.809017
			y: 2.118034
			z: 1.0
		}, Vertex{
			x: -0.809017
			y: 2.118034
			z: -1.0
		}, Vertex{
			x: -0.809017
			y: -2.118034
			z: 1.0
		}, Vertex{
			x: -0.809017
			y: -2.118034
			z: -1.0
		}, Vertex{
			x: 0.5
			y: 1.618034
			z: 1.809017
		}, Vertex{
			x: 0.5
			y: 1.618034
			z: -1.809017
		}, Vertex{
			x: 0.5
			y: -1.618034
			z: 1.809017
		}, Vertex{
			x: 0.5
			y: -1.618034
			z: -1.809017
		}, Vertex{
			x: -0.5
			y: 1.618034
			z: 1.809017
		}, Vertex{
			x: -0.5
			y: 1.618034
			z: -1.809017
		}, Vertex{
			x: -0.5
			y: -1.618034
			z: 1.809017
		}, Vertex{
			x: -0.5
			y: -1.618034
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.5
			z: 1.618034
		}, Vertex{
			x: 1.809017
			y: 0.5
			z: -1.618034
		}, Vertex{
			x: 1.809017
			y: -0.5
			z: 1.618034
		}, Vertex{
			x: 1.809017
			y: -0.5
			z: -1.618034
		}, Vertex{
			x: -1.809017
			y: 0.5
			z: 1.618034
		}, Vertex{
			x: -1.809017
			y: 0.5
			z: -1.618034
		}, Vertex{
			x: -1.809017
			y: -0.5
			z: 1.618034
		}, Vertex{
			x: -1.809017
			y: -0.5
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 1.809017
			z: 0.5
		}, Vertex{
			x: 1.618034
			y: 1.809017
			z: -0.5
		}, Vertex{
			x: 1.618034
			y: -1.809017
			z: 0.5
		}, Vertex{
			x: 1.618034
			y: -1.809017
			z: -0.5
		}, Vertex{
			x: -1.618034
			y: 1.809017
			z: 0.5
		}, Vertex{
			x: -1.618034
			y: 1.809017
			z: -0.5
		}, Vertex{
			x: -1.618034
			y: -1.809017
			z: 0.5
		}, Vertex{
			x: -1.618034
			y: -1.809017
			z: -0.5
		}]
		faces:     [[0, 2, 18, 42, 38, 14], [1, 3, 17, 41, 37, 13],
			[2, 0, 12, 36, 40, 16], [3, 1, 15, 39, 43, 19], [4, 5, 23, 47, 45, 21],
			[5, 4, 20, 44, 46, 22], [6, 7, 26, 50, 48, 24], [7, 6, 25, 49, 51, 27],
			[8, 9, 33, 57, 56, 32], [9, 8, 28, 52, 53, 29], [10, 11, 31, 55, 54, 30],
			[11, 10, 34, 58, 59, 35], [12, 44, 20, 52, 28, 36],
			[13, 37, 29, 53, 21, 45], [14, 38, 30, 54, 22, 46],
			[15, 47, 23, 55, 31, 39], [16, 40, 32, 56, 24, 48],
			[17, 49, 25, 57, 33, 41], [18, 50, 26, 58, 34, 42],
			[19, 43, 35, 59, 27, 51], [0, 14, 46, 44, 12], [1, 13, 45, 47, 15],
			[2, 16, 48, 50, 18], [3, 19, 51, 49, 17], [4, 21, 53, 52, 20],
			[5, 22, 54, 55, 23], [6, 24, 56, 57, 25], [7, 27, 59, 58, 26],
			[8, 32, 40, 36, 28], [9, 29, 37, 41, 33], [10, 30, 38, 42, 34],
			[11, 35, 43, 39, 31]]
	},
	Polyhedron{
		name:      'Octahemioctahedron'
		vertexes_: [Vertex{
			x: 0.7071068
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: 0.7071068
		}, Vertex{
			x: -0.7071068
			y: 0.0
			z: -0.7071068
		}, Vertex{
			x: 0.7071068
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: 0.7071068
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: 0.7071068
			z: 0.0
		}, Vertex{
			x: -0.7071068
			y: -0.7071068
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: 0.7071068
			z: -0.7071068
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: 0.7071068
		}, Vertex{
			x: 0.0
			y: -0.7071068
			z: -0.7071068
		}]
		faces:     [[0, 4, 9, 3, 7, 10], [0, 5, 11, 3, 6, 8],
			[1, 4, 8, 2, 7, 11], [1, 5, 10, 2, 6, 9], [0, 8, 4],
			[0, 10, 5], [1, 9, 4], [1, 11, 5], [2, 8, 6], [2, 10, 7],
			[3, 9, 6], [3, 11, 7]]
	},
	Polyhedron{
		name:      'GreatSnubDodecicosidodecahedron'
		vertexes_: [Vertex{
			x: 0.1817730
			y: 0.1429011
			z: 0.6682349
		}, Vertex{
			x: 0.1817730
			y: 0.1429011
			z: -0.6682349
		}, Vertex{
			x: 0.1817730
			y: -0.1429011
			z: 0.6682349
		}, Vertex{
			x: 0.1817730
			y: -0.1429011
			z: -0.6682349
		}, Vertex{
			x: -0.1817730
			y: 0.1429011
			z: 0.6682349
		}, Vertex{
			x: -0.1817730
			y: 0.1429011
			z: -0.6682349
		}, Vertex{
			x: -0.1817730
			y: -0.1429011
			z: 0.6682349
		}, Vertex{
			x: -0.1817730
			y: -0.1429011
			z: -0.6682349
		}, Vertex{
			x: 0.6682349
			y: 0.1817730
			z: 0.1429011
		}, Vertex{
			x: 0.6682349
			y: 0.1817730
			z: -0.1429011
		}, Vertex{
			x: 0.6682349
			y: -0.1817730
			z: 0.1429011
		}, Vertex{
			x: 0.6682349
			y: -0.1817730
			z: -0.1429011
		}, Vertex{
			x: -0.6682349
			y: 0.1817730
			z: 0.1429011
		}, Vertex{
			x: -0.6682349
			y: 0.1817730
			z: -0.1429011
		}, Vertex{
			x: -0.6682349
			y: -0.1817730
			z: 0.1429011
		}, Vertex{
			x: -0.6682349
			y: -0.1817730
			z: -0.1429011
		}, Vertex{
			x: 0.1429011
			y: 0.6682349
			z: 0.1817730
		}, Vertex{
			x: 0.1429011
			y: 0.6682349
			z: -0.1817730
		}, Vertex{
			x: 0.1429011
			y: -0.6682349
			z: 0.1817730
		}, Vertex{
			x: 0.1429011
			y: -0.6682349
			z: -0.1817730
		}, Vertex{
			x: -0.1429011
			y: 0.6682349
			z: 0.1817730
		}, Vertex{
			x: -0.1429011
			y: 0.6682349
			z: -0.1817730
		}, Vertex{
			x: -0.1429011
			y: -0.6682349
			z: 0.1817730
		}, Vertex{
			x: -0.1429011
			y: -0.6682349
			z: -0.1817730
		}, Vertex{
			x: 0.0
			y: 0.437016
			z: 0.5558929
		}, Vertex{
			x: 0.0
			y: 0.437016
			z: -0.5558929
		}, Vertex{
			x: 0.0
			y: -0.437016
			z: 0.5558929
		}, Vertex{
			x: 0.0
			y: -0.437016
			z: -0.5558929
		}, Vertex{
			x: 0.5558929
			y: 0.0
			z: 0.437016
		}, Vertex{
			x: 0.5558929
			y: 0.0
			z: -0.437016
		}, Vertex{
			x: -0.5558929
			y: 0.0
			z: 0.437016
		}, Vertex{
			x: -0.5558929
			y: 0.0
			z: -0.437016
		}, Vertex{
			x: 0.437016
			y: 0.5558929
			z: 0.0
		}, Vertex{
			x: 0.437016
			y: -0.5558929
			z: 0.0
		}, Vertex{
			x: -0.437016
			y: 0.5558929
			z: 0.0
		}, Vertex{
			x: -0.437016
			y: -0.5558929
			z: 0.0
		}, Vertex{
			x: 0.4129919
			y: 0.2312188
			z: 0.5253338
		}, Vertex{
			x: 0.4129919
			y: 0.2312188
			z: -0.5253338
		}, Vertex{
			x: 0.4129919
			y: -0.2312188
			z: 0.5253338
		}, Vertex{
			x: 0.4129919
			y: -0.2312188
			z: -0.5253338
		}, Vertex{
			x: -0.4129919
			y: 0.2312188
			z: 0.5253338
		}, Vertex{
			x: -0.4129919
			y: 0.2312188
			z: -0.5253338
		}, Vertex{
			x: -0.4129919
			y: -0.2312188
			z: 0.5253338
		}, Vertex{
			x: -0.4129919
			y: -0.2312188
			z: -0.5253338
		}, Vertex{
			x: 0.5253338
			y: 0.4129919
			z: 0.2312188
		}, Vertex{
			x: 0.5253338
			y: 0.4129919
			z: -0.2312188
		}, Vertex{
			x: 0.5253338
			y: -0.4129919
			z: 0.2312188
		}, Vertex{
			x: 0.5253338
			y: -0.4129919
			z: -0.2312188
		}, Vertex{
			x: -0.5253338
			y: 0.4129919
			z: 0.2312188
		}, Vertex{
			x: -0.5253338
			y: 0.4129919
			z: -0.2312188
		}, Vertex{
			x: -0.5253338
			y: -0.4129919
			z: 0.2312188
		}, Vertex{
			x: -0.5253338
			y: -0.4129919
			z: -0.2312188
		}, Vertex{
			x: 0.2312188
			y: 0.5253338
			z: 0.4129919
		}, Vertex{
			x: 0.2312188
			y: 0.5253338
			z: -0.4129919
		}, Vertex{
			x: 0.2312188
			y: -0.5253338
			z: 0.4129919
		}, Vertex{
			x: 0.2312188
			y: -0.5253338
			z: -0.4129919
		}, Vertex{
			x: -0.2312188
			y: 0.5253338
			z: 0.4129919
		}, Vertex{
			x: -0.2312188
			y: 0.5253338
			z: -0.4129919
		}, Vertex{
			x: -0.2312188
			y: -0.5253338
			z: 0.4129919
		}, Vertex{
			x: -0.2312188
			y: -0.5253338
			z: -0.4129919
		}]
		faces:     [[16, 10, 53, 36, 29], [16, 41, 45, 34, 1],
			[17, 11, 52, 37, 28], [17, 40, 44, 34, 0], [18, 8, 55, 38, 29],
			[18, 43, 47, 35, 3], [19, 9, 54, 39, 28], [19, 42, 46, 35, 2],
			[20, 14, 57, 40, 31], [20, 37, 49, 32, 5], [21, 15, 56, 41, 30],
			[21, 36, 48, 32, 4], [22, 12, 59, 42, 31], [22, 39, 51, 33, 7],
			[23, 13, 58, 43, 30], [23, 38, 50, 33, 6], [24, 10, 6, 44, 54],
			[24, 14, 2, 48, 58], [25, 11, 7, 45, 55], [25, 15, 3, 49, 59],
			[26, 8, 4, 46, 52], [26, 12, 0, 50, 56], [27, 9, 5, 47, 53],
			[27, 13, 1, 51, 57], [0, 34, 50], [1, 13, 16], [2, 14, 19],
			[3, 35, 49], [4, 8, 21], [5, 32, 47], [6, 33, 44],
			[7, 11, 22], [8, 26, 55], [9, 19, 5], [10, 16, 6],
			[11, 25, 52], [12, 22, 0], [13, 27, 58], [14, 24, 57],
			[15, 21, 3], [16, 29, 41], [17, 0, 11], [18, 3, 8],
			[19, 28, 42], [20, 5, 14], [21, 30, 36], [22, 31, 39],
			[23, 6, 13], [24, 58, 10], [25, 55, 15], [26, 52, 12],
			[27, 57, 9], [28, 39, 17], [29, 36, 18], [30, 41, 23],
			[31, 42, 20], [32, 49, 4], [33, 50, 7], [34, 44, 1],
			[35, 47, 2], [36, 53, 48], [37, 20, 28], [38, 23, 29],
			[39, 54, 51], [40, 17, 31], [41, 56, 45], [42, 59, 46],
			[43, 18, 30], [44, 40, 54], [45, 7, 34], [46, 4, 35],
			[47, 43, 53], [48, 2, 32], [49, 37, 59], [50, 38, 56],
			[51, 1, 33], [52, 46, 37], [53, 10, 27], [54, 9, 24],
			[55, 45, 38], [56, 15, 26], [57, 51, 40], [58, 48, 43],
			[59, 12, 25], [0, 22, 11], [1, 44, 33], [2, 47, 32],
			[3, 21, 8], [4, 49, 35], [5, 19, 14], [6, 16, 13],
			[7, 50, 34], [28, 20, 42], [29, 23, 41], [30, 18, 36],
			[31, 17, 39], [52, 25, 12], [53, 43, 48], [54, 40, 51],
			[55, 26, 15], [56, 38, 45], [57, 24, 9], [58, 27, 10],
			[59, 37, 46]]
	},
	Polyhedron{
		name:      'TruncatedTetrahedron'
		vertexes_: [Vertex{
			x: 0.3535534
			y: -0.3535534
			z: 1.060660
		}, Vertex{
			x: 0.3535534
			y: 0.3535534
			z: -1.060660
		}, Vertex{
			x: -0.3535534
			y: 0.3535534
			z: 1.060660
		}, Vertex{
			x: -0.3535534
			y: -0.3535534
			z: -1.060660
		}, Vertex{
			x: 1.060660
			y: -0.3535534
			z: 0.3535534
		}, Vertex{
			x: 1.060660
			y: 0.3535534
			z: -0.3535534
		}, Vertex{
			x: -1.060660
			y: 0.3535534
			z: 0.3535534
		}, Vertex{
			x: -1.060660
			y: -0.3535534
			z: -0.3535534
		}, Vertex{
			x: 0.3535534
			y: -1.060660
			z: 0.3535534
		}, Vertex{
			x: 0.3535534
			y: 1.060660
			z: -0.3535534
		}, Vertex{
			x: -0.3535534
			y: 1.060660
			z: 0.3535534
		}, Vertex{
			x: -0.3535534
			y: -1.060660
			z: -0.3535534
		}]
		faces:     [[0, 4, 5, 9, 10, 2], [1, 5, 4, 8, 11, 3],
			[2, 6, 7, 11, 8, 0], [3, 7, 6, 10, 9, 1], [0, 8, 4],
			[1, 9, 5], [2, 10, 6], [3, 11, 7]]
	},
	Polyhedron{
		name:      'SmallDodecahemicosahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: -0.309017
		}, Vertex{
			x: 0.809017
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: -0.809017
		}]
		faces:     [[0, 14, 15, 1, 21, 20], [0, 16, 17, 1, 19, 18],
			[2, 22, 26, 3, 29, 25], [2, 23, 27, 3, 28, 24], [4, 6, 8, 5, 13, 11],
			[4, 7, 9, 5, 12, 10], [6, 16, 25, 13, 19, 26], [7, 17, 24, 12, 18, 27],
			[8, 14, 23, 11, 21, 28], [9, 15, 22, 10, 20, 29],
			[0, 14, 23, 27, 18], [0, 20, 29, 25, 16], [1, 17, 24, 28, 21],
			[1, 19, 26, 22, 15], [2, 22, 10, 12, 24], [2, 25, 13, 11, 23],
			[3, 27, 7, 9, 29], [3, 28, 8, 6, 26], [4, 6, 16, 17, 7],
			[4, 11, 21, 20, 10], [5, 12, 18, 19, 13], [5, 9, 15, 14, 8]]
	},
	Polyhedron{
		name:      'GreatDodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.0
			z: 0.809017
		}, Vertex{
			x: 0.5
			y: 0.0
			z: -0.809017
		}, Vertex{
			x: -0.5
			y: 0.0
			z: 0.809017
		}, Vertex{
			x: -0.5
			y: 0.0
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.5
			z: 0.0
		}, Vertex{
			x: 0.809017
			y: -0.5
			z: 0.0
		}, Vertex{
			x: -0.809017
			y: 0.5
			z: 0.0
		}, Vertex{
			x: -0.809017
			y: -0.5
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.809017
			z: 0.5
		}, Vertex{
			x: 0.0
			y: 0.809017
			z: -0.5
		}, Vertex{
			x: 0.0
			y: -0.809017
			z: 0.5
		}, Vertex{
			x: 0.0
			y: -0.809017
			z: -0.5
		}]
		faces:     [[0, 2, 7, 11, 5], [0, 5, 1, 9, 8], [0, 8, 6, 7, 10],
			[1, 3, 6, 8, 4], [1, 4, 0, 10, 11], [1, 11, 7, 6, 9],
			[2, 0, 4, 9, 6], [2, 6, 3, 11, 10], [2, 10, 5, 4, 8],
			[3, 1, 5, 10, 7], [3, 7, 2, 8, 9], [3, 9, 4, 5, 11]]
	},
	Polyhedron{
		name:      'GreatTriakisIcosahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.690983
			z: -0.4270510
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -0.4270510
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.690983
			y: -0.4270510
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -0.4270510
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: 0.4270510
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 0.4270510
			z: 0.0
		}, Vertex{
			x: -0.4270510
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -0.4270510
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.4270510
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.4270510
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.5413559
			y: 0.0
			z: 0.2067796
		}, Vertex{
			x: 0.5413559
			y: 0.0
			z: -0.2067796
		}, Vertex{
			x: -0.5413559
			y: 0.0
			z: 0.2067796
		}, Vertex{
			x: -0.5413559
			y: 0.0
			z: -0.2067796
		}, Vertex{
			x: 0.0
			y: 0.2067796
			z: 0.5413559
		}, Vertex{
			x: 0.0
			y: 0.2067796
			z: -0.5413559
		}, Vertex{
			x: 0.0
			y: -0.2067796
			z: 0.5413559
		}, Vertex{
			x: 0.0
			y: -0.2067796
			z: -0.5413559
		}, Vertex{
			x: 0.2067796
			y: 0.5413559
			z: 0.0
		}, Vertex{
			x: -0.2067796
			y: 0.5413559
			z: 0.0
		}, Vertex{
			x: 0.2067796
			y: -0.5413559
			z: 0.0
		}, Vertex{
			x: -0.2067796
			y: -0.5413559
			z: 0.0
		}, Vertex{
			x: -0.3345763
			y: -0.3345763
			z: -0.3345763
		}, Vertex{
			x: -0.3345763
			y: -0.3345763
			z: 0.3345763
		}, Vertex{
			x: 0.3345763
			y: -0.3345763
			z: -0.3345763
		}, Vertex{
			x: 0.3345763
			y: -0.3345763
			z: 0.3345763
		}, Vertex{
			x: -0.3345763
			y: 0.3345763
			z: -0.3345763
		}, Vertex{
			x: -0.3345763
			y: 0.3345763
			z: 0.3345763
		}, Vertex{
			x: 0.3345763
			y: 0.3345763
			z: -0.3345763
		}, Vertex{
			x: 0.3345763
			y: 0.3345763
			z: 0.3345763
		}]
		faces:     [[12, 0, 8], [12, 8, 2], [12, 2, 0], [13, 1, 3],
			[13, 3, 9], [13, 9, 1], [14, 0, 2], [14, 2, 10], [14, 10, 0],
			[15, 1, 11], [15, 11, 3], [15, 3, 1], [16, 0, 5],
			[16, 5, 4], [16, 4, 0], [17, 1, 4], [17, 4, 5], [17, 5, 1],
			[18, 2, 6], [18, 6, 7], [18, 7, 2], [19, 3, 7], [19, 7, 6],
			[19, 6, 3], [20, 4, 9], [20, 9, 8], [20, 8, 4], [21, 5, 10],
			[21, 10, 11], [21, 11, 5], [22, 6, 8], [22, 8, 9],
			[22, 9, 6], [23, 7, 11], [23, 11, 10], [23, 10, 7],
			[24, 0, 4], [24, 4, 8], [24, 8, 0], [25, 1, 9], [25, 9, 4],
			[25, 4, 1], [26, 0, 10], [26, 10, 5], [26, 5, 0],
			[27, 1, 5], [27, 5, 11], [27, 11, 1], [28, 2, 8],
			[28, 8, 6], [28, 6, 2], [29, 3, 6], [29, 6, 9], [29, 9, 3],
			[30, 2, 7], [30, 7, 10], [30, 10, 2], [31, 3, 11],
			[31, 11, 7], [31, 7, 3]]
	},
	Polyhedron{
		name:      'SnubDodecahedron(dextro}'
		vertexes_: [Vertex{
			x: 0.3748217
			y: 0.3309210
			z: 2.097054
		}, Vertex{
			x: 0.3748217
			y: -0.3309210
			z: -2.097054
		}, Vertex{
			x: -0.3748217
			y: -0.3309210
			z: 2.097054
		}, Vertex{
			x: -0.3748217
			y: 0.3309210
			z: -2.097054
		}, Vertex{
			x: 2.097054
			y: 0.3748217
			z: 0.3309210
		}, Vertex{
			x: 2.097054
			y: -0.3748217
			z: -0.3309210
		}, Vertex{
			x: -2.097054
			y: -0.3748217
			z: 0.3309210
		}, Vertex{
			x: -2.097054
			y: 0.3748217
			z: -0.3309210
		}, Vertex{
			x: 0.3309210
			y: 2.097054
			z: 0.3748217
		}, Vertex{
			x: 0.3309210
			y: -2.097054
			z: -0.3748217
		}, Vertex{
			x: -0.3309210
			y: -2.097054
			z: 0.3748217
		}, Vertex{
			x: -0.3309210
			y: 2.097054
			z: -0.3748217
		}, Vertex{
			x: 0.5677154
			y: -0.6430296
			z: 1.977839
		}, Vertex{
			x: 0.5677154
			y: 0.6430296
			z: -1.977839
		}, Vertex{
			x: -0.5677154
			y: 0.6430296
			z: 1.977839
		}, Vertex{
			x: -0.5677154
			y: -0.6430296
			z: -1.977839
		}, Vertex{
			x: 1.977839
			y: -0.5677154
			z: 0.6430296
		}, Vertex{
			x: 1.977839
			y: 0.5677154
			z: -0.6430296
		}, Vertex{
			x: -1.977839
			y: 0.5677154
			z: 0.6430296
		}, Vertex{
			x: -1.977839
			y: -0.5677154
			z: -0.6430296
		}, Vertex{
			x: 0.6430296
			y: -1.977839
			z: 0.5677154
		}, Vertex{
			x: 0.6430296
			y: 1.977839
			z: -0.5677154
		}, Vertex{
			x: -0.6430296
			y: 1.977839
			z: 0.5677154
		}, Vertex{
			x: -0.6430296
			y: -1.977839
			z: -0.5677154
		}, Vertex{
			x: 0.1928937
			y: 1.249504
			z: 1.746187
		}, Vertex{
			x: 0.1928937
			y: -1.249504
			z: -1.746187
		}, Vertex{
			x: -0.1928937
			y: -1.249504
			z: 1.746187
		}, Vertex{
			x: -0.1928937
			y: 1.249504
			z: -1.746187
		}, Vertex{
			x: 1.746187
			y: 0.1928937
			z: 1.249504
		}, Vertex{
			x: 1.746187
			y: -0.1928937
			z: -1.249504
		}, Vertex{
			x: -1.746187
			y: -0.1928937
			z: 1.249504
		}, Vertex{
			x: -1.746187
			y: 0.1928937
			z: -1.249504
		}, Vertex{
			x: 1.249504
			y: 1.746187
			z: 0.1928937
		}, Vertex{
			x: 1.249504
			y: -1.746187
			z: -0.1928937
		}, Vertex{
			x: -1.249504
			y: -1.746187
			z: 0.1928937
		}, Vertex{
			x: -1.249504
			y: 1.746187
			z: -0.1928937
		}, Vertex{
			x: 1.103157
			y: 0.8475500
			z: 1.646918
		}, Vertex{
			x: 1.103157
			y: -0.8475500
			z: -1.646918
		}, Vertex{
			x: -1.103157
			y: -0.8475500
			z: 1.646918
		}, Vertex{
			x: -1.103157
			y: 0.8475500
			z: -1.646918
		}, Vertex{
			x: 1.646918
			y: 1.103157
			z: 0.8475500
		}, Vertex{
			x: 1.646918
			y: -1.103157
			z: -0.8475500
		}, Vertex{
			x: -1.646918
			y: -1.103157
			z: 0.8475500
		}, Vertex{
			x: -1.646918
			y: 1.103157
			z: -0.8475500
		}, Vertex{
			x: 0.8475500
			y: 1.646918
			z: 1.103157
		}, Vertex{
			x: 0.8475500
			y: -1.646918
			z: -1.103157
		}, Vertex{
			x: -0.8475500
			y: -1.646918
			z: 1.103157
		}, Vertex{
			x: -0.8475500
			y: 1.646918
			z: -1.103157
		}, Vertex{
			x: 1.415265
			y: -0.7283352
			z: 1.454024
		}, Vertex{
			x: 1.415265
			y: 0.7283352
			z: -1.454024
		}, Vertex{
			x: -1.415265
			y: 0.7283352
			z: 1.454024
		}, Vertex{
			x: -1.415265
			y: -0.7283352
			z: -1.454024
		}, Vertex{
			x: 1.454024
			y: -1.415265
			z: 0.7283352
		}, Vertex{
			x: 1.454024
			y: 1.415265
			z: -0.7283352
		}, Vertex{
			x: -1.454024
			y: 1.415265
			z: 0.7283352
		}, Vertex{
			x: -1.454024
			y: -1.415265
			z: -0.7283352
		}, Vertex{
			x: 0.7283352
			y: -1.454024
			z: 1.415265
		}, Vertex{
			x: 0.7283352
			y: 1.454024
			z: -1.415265
		}, Vertex{
			x: -0.7283352
			y: 1.454024
			z: 1.415265
		}, Vertex{
			x: -0.7283352
			y: -1.454024
			z: -1.415265
		}]
		faces:     [[0, 12, 48, 28, 36], [1, 13, 49, 29, 37],
			[2, 14, 50, 30, 38], [3, 15, 51, 31, 39], [4, 17, 53, 32, 40],
			[5, 16, 52, 33, 41], [6, 19, 55, 34, 42], [7, 18, 54, 35, 43],
			[8, 22, 58, 24, 44], [9, 23, 59, 25, 45], [10, 20, 56, 26, 46],
			[11, 21, 57, 27, 47], [0, 14, 2], [1, 15, 3], [2, 12, 0],
			[3, 13, 1], [4, 16, 5], [5, 17, 4], [6, 18, 7], [7, 19, 6],
			[8, 21, 11], [9, 20, 10], [10, 23, 9], [11, 22, 8],
			[12, 56, 48], [13, 57, 49], [14, 58, 50], [15, 59, 51],
			[16, 48, 52], [17, 49, 53], [18, 50, 54], [19, 51, 55],
			[20, 52, 56], [21, 53, 57], [22, 54, 58], [23, 55, 59],
			[24, 36, 44], [25, 37, 45], [26, 38, 46], [27, 39, 47],
			[28, 40, 36], [29, 41, 37], [30, 42, 38], [31, 43, 39],
			[32, 44, 40], [33, 45, 41], [34, 46, 42], [35, 47, 43],
			[36, 24, 0], [37, 25, 1], [38, 26, 2], [39, 27, 3],
			[40, 28, 4], [41, 29, 5], [42, 30, 6], [43, 31, 7],
			[44, 32, 8], [45, 33, 9], [46, 34, 10], [47, 35, 11],
			[48, 16, 28], [49, 17, 29], [50, 18, 30], [51, 19, 31],
			[52, 20, 33], [53, 21, 32], [54, 22, 35], [55, 23, 34],
			[56, 12, 26], [57, 13, 27], [58, 14, 24], [59, 15, 25],
			[24, 14, 0], [25, 15, 1], [26, 12, 2], [27, 13, 3],
			[28, 16, 4], [29, 17, 5], [30, 18, 6], [31, 19, 7],
			[32, 21, 8], [33, 20, 9], [34, 23, 10], [35, 22, 11],
			[36, 40, 44], [37, 41, 45], [38, 42, 46], [39, 43, 47],
			[48, 56, 52], [49, 57, 53], [50, 58, 54], [51, 59, 55]]
	},
	Polyhedron{
		name:      'TetrakisHexahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.590990
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.590990
		}, Vertex{
			x: 1.590990
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.590990
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.590990
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.590990
			z: 0.0
		}, Vertex{
			x: 1.060660
			y: 1.060660
			z: 1.060660
		}, Vertex{
			x: 1.060660
			y: 1.060660
			z: -1.060660
		}, Vertex{
			x: 1.060660
			y: -1.060660
			z: 1.060660
		}, Vertex{
			x: 1.060660
			y: -1.060660
			z: -1.060660
		}, Vertex{
			x: -1.060660
			y: 1.060660
			z: 1.060660
		}, Vertex{
			x: -1.060660
			y: 1.060660
			z: -1.060660
		}, Vertex{
			x: -1.060660
			y: -1.060660
			z: 1.060660
		}, Vertex{
			x: -1.060660
			y: -1.060660
			z: -1.060660
		}]
		faces:     [[0, 6, 10], [0, 10, 12], [0, 12, 8], [0, 8, 6],
			[1, 7, 9], [1, 9, 13], [1, 13, 11], [1, 11, 7], [2, 6, 8],
			[2, 8, 9], [2, 9, 7], [2, 7, 6], [3, 10, 11], [3, 11, 13],
			[3, 13, 12], [3, 12, 10], [4, 6, 7], [4, 7, 11], [4, 11, 10],
			[4, 10, 6], [5, 8, 12], [5, 12, 13], [5, 13, 9], [5, 9, 8]]
	},
	Polyhedron{
		name:      'TruncatedCube'
		vertexes_: [Vertex{
			x: 1.207107
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: 1.207107
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: 1.207107
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: 1.207107
		}, Vertex{
			x: -1.207107
			y: 0.5
			z: -1.207107
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: 1.207107
		}, Vertex{
			x: -1.207107
			y: -0.5
			z: -1.207107
		}, Vertex{
			x: 1.207107
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: 1.207107
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: 1.207107
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: 1.207107
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: 1.207107
			z: -0.5
		}, Vertex{
			x: -1.207107
			y: -1.207107
			z: 0.5
		}, Vertex{
			x: -1.207107
			y: -1.207107
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: 1.207107
			z: -1.207107
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: 1.207107
		}, Vertex{
			x: 0.5
			y: -1.207107
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: 1.207107
			z: -1.207107
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: 1.207107
		}, Vertex{
			x: -0.5
			y: -1.207107
			z: -1.207107
		}]
		faces:     [[0, 2, 10, 11, 3, 1, 9, 8], [0, 16, 20, 4, 6, 22, 18, 2],
			[12, 13, 5, 7, 15, 14, 6, 4], [12, 20, 16, 8, 9, 17, 21, 13],
			[19, 23, 7, 5, 21, 17, 1, 3], [19, 11, 10, 18, 22, 14, 15, 23],
			[0, 8, 16], [1, 17, 9], [2, 18, 10], [3, 11, 19],
			[4, 20, 12], [5, 13, 21], [6, 14, 22], [7, 23, 15]]
	},
	Polyhedron{
		name:      'GreatDisdyakisDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.9611318
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.9611318
		}, Vertex{
			x: 0.9611318
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.9611318
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.9611318
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.9611318
			z: 0.0
		}, Vertex{
			x: 0.7836116
			y: 0.0
			z: 0.7836116
		}, Vertex{
			x: 0.7836116
			y: 0.0
			z: -0.7836116
		}, Vertex{
			x: -0.7836116
			y: 0.0
			z: 0.7836116
		}, Vertex{
			x: -0.7836116
			y: 0.0
			z: -0.7836116
		}, Vertex{
			x: 0.7836116
			y: 0.7836116
			z: 0.0
		}, Vertex{
			x: 0.7836116
			y: -0.7836116
			z: 0.0
		}, Vertex{
			x: -0.7836116
			y: 0.7836116
			z: 0.0
		}, Vertex{
			x: -0.7836116
			y: -0.7836116
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.7836116
			z: 0.7836116
		}, Vertex{
			x: 0.0
			y: 0.7836116
			z: -0.7836116
		}, Vertex{
			x: 0.0
			y: -0.7836116
			z: 0.7836116
		}, Vertex{
			x: 0.0
			y: -0.7836116
			z: -0.7836116
		}, Vertex{
			x: 1.414214
			y: 1.414214
			z: 1.414214
		}, Vertex{
			x: 1.414214
			y: 1.414214
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: -1.414214
			z: 1.414214
		}, Vertex{
			x: 1.414214
			y: -1.414214
			z: -1.414214
		}, Vertex{
			x: -1.414214
			y: 1.414214
			z: 1.414214
		}, Vertex{
			x: -1.414214
			y: 1.414214
			z: -1.414214
		}, Vertex{
			x: -1.414214
			y: -1.414214
			z: 1.414214
		}, Vertex{
			x: -1.414214
			y: -1.414214
			z: -1.414214
		}]
		faces:     [[0, 6, 18], [0, 18, 14], [0, 14, 22], [0, 22, 8],
			[0, 8, 24], [0, 24, 16], [0, 16, 20], [0, 20, 6],
			[1, 7, 21], [1, 21, 17], [1, 17, 25], [1, 25, 9],
			[1, 9, 23], [1, 23, 15], [1, 15, 19], [1, 19, 7],
			[2, 6, 20], [2, 20, 11], [2, 11, 21], [2, 21, 7],
			[2, 7, 19], [2, 19, 10], [2, 10, 18], [2, 18, 6],
			[3, 8, 22], [3, 22, 12], [3, 12, 23], [3, 23, 9],
			[3, 9, 25], [3, 25, 13], [3, 13, 24], [3, 24, 8],
			[4, 10, 19], [4, 19, 15], [4, 15, 23], [4, 23, 12],
			[4, 12, 22], [4, 22, 14], [4, 14, 18], [4, 18, 10],
			[5, 11, 20], [5, 20, 16], [5, 16, 24], [5, 24, 13],
			[5, 13, 25], [5, 25, 17], [5, 17, 21], [5, 21, 11]]
	},
	Polyhedron{
		name:      'GreatPentakisDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.690983
			z: -0.4270510
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -0.4270510
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.690983
			y: -0.4270510
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -0.4270510
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: 0.4270510
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 0.4270510
			z: 0.0
		}, Vertex{
			x: -0.4270510
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -0.4270510
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.4270510
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.4270510
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.0
			y: 6.545085
			z: -4.045085
		}, Vertex{
			x: 0.0
			y: 6.545085
			z: 4.045085
		}, Vertex{
			x: 0.0
			y: -6.545085
			z: -4.045085
		}, Vertex{
			x: 0.0
			y: -6.545085
			z: 4.045085
		}, Vertex{
			x: 6.545085
			y: -4.045085
			z: 0.0
		}, Vertex{
			x: -6.545085
			y: -4.045085
			z: 0.0
		}, Vertex{
			x: 6.545085
			y: 4.045085
			z: 0.0
		}, Vertex{
			x: -6.545085
			y: 4.045085
			z: 0.0
		}, Vertex{
			x: -4.045085
			y: 0.0
			z: 6.545085
		}, Vertex{
			x: -4.045085
			y: 0.0
			z: -6.545085
		}, Vertex{
			x: 4.045085
			y: 0.0
			z: 6.545085
		}, Vertex{
			x: 4.045085
			y: 0.0
			z: -6.545085
		}]
		faces:     [[12, 2, 5], [12, 5, 8], [12, 8, 10], [12, 10, 4],
			[12, 4, 2], [13, 3, 4], [13, 4, 11], [13, 11, 9],
			[13, 9, 5], [13, 5, 3], [14, 0, 6], [14, 6, 10], [14, 10, 8],
			[14, 8, 7], [14, 7, 0], [15, 1, 7], [15, 7, 9], [15, 9, 11],
			[15, 11, 6], [15, 6, 1], [16, 0, 1], [16, 1, 8], [16, 8, 5],
			[16, 5, 9], [16, 9, 0], [17, 1, 0], [17, 0, 11], [17, 11, 4],
			[17, 4, 10], [17, 10, 1], [18, 3, 2], [18, 2, 9],
			[18, 9, 7], [18, 7, 8], [18, 8, 3], [19, 2, 3], [19, 3, 10],
			[19, 10, 6], [19, 6, 11], [19, 11, 2], [20, 0, 9],
			[20, 9, 2], [20, 2, 4], [20, 4, 6], [20, 6, 0], [21, 1, 6],
			[21, 6, 4], [21, 4, 3], [21, 3, 8], [21, 8, 1], [22, 0, 7],
			[22, 7, 5], [22, 5, 2], [22, 2, 11], [22, 11, 0],
			[23, 1, 10], [23, 10, 3], [23, 3, 5], [23, 5, 7],
			[23, 7, 1]]
	},
	Polyhedron{
		name:      'MedialTriambicIcosahedron'
		vertexes_: [Vertex{
			x: 1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: 1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: 2.618034
		}, Vertex{
			x: -1.618034
			y: 0.0
			z: -2.618034
		}, Vertex{
			x: 2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: 2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: 1.618034
			z: 0.0
		}, Vertex{
			x: -2.618034
			y: -1.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: 2.618034
			z: -1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: 1.618034
		}, Vertex{
			x: 0.0
			y: -2.618034
			z: -1.618034
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: -0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: -0.3819660
		}]
		faces:     [[0, 14, 6, 19, 11, 22], [0, 22, 7, 23, 1, 17],
			[0, 17, 11, 13, 9, 16], [0, 16, 1, 21, 6, 20], [0, 20, 9, 18, 7, 14],
			[3, 13, 4, 17, 10, 23], [3, 23, 5, 22, 2, 19], [3, 19, 10, 14, 8, 18],
			[3, 18, 2, 20, 4, 21], [3, 21, 8, 16, 5, 13], [12, 2, 22, 11, 17, 4],
			[12, 4, 20, 6, 14, 10], [12, 10, 17, 1, 16, 8], [12, 8, 14, 7, 22, 5],
			[12, 5, 16, 9, 20, 2], [15, 1, 23, 10, 19, 6], [15, 6, 21, 4, 13, 11],
			[15, 11, 19, 2, 18, 9], [15, 9, 13, 5, 23, 7], [15, 7, 18, 8, 21, 1]]
	},
	Polyhedron{
		name:      'SmallStellatedTruncatedDodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.5
			z: 0.690983
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -0.690983
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 0.690983
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -0.690983
		}, Vertex{
			x: 0.5
			y: 0.690983
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 0.690983
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -0.690983
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -0.690983
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 0.690983
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -0.690983
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -0.690983
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: -0.618034
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: 0.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: -0.618034
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: 0.618034
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: -0.618034
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: 0.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: -0.618034
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: 0.618034
		}, Vertex{
			x: -0.309017
			y: -0.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: -0.618034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: -0.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: -0.618034
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: 0.618034
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: 0.618034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 0.618034
			z: 0.5
		}, Vertex{
			x: 0.309017
			y: 0.618034
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: -0.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: 0.618034
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: 0.618034
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: -0.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: -0.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 0.618034
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: 0.618034
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: 0.1909830
			z: 0.1909830
		}, Vertex{
			x: -0.809017
			y: 0.1909830
			z: -0.1909830
		}, Vertex{
			x: 0.809017
			y: 0.1909830
			z: 0.1909830
		}, Vertex{
			x: 0.809017
			y: 0.1909830
			z: -0.1909830
		}, Vertex{
			x: -0.809017
			y: -0.1909830
			z: 0.1909830
		}, Vertex{
			x: -0.809017
			y: -0.1909830
			z: -0.1909830
		}, Vertex{
			x: 0.809017
			y: -0.1909830
			z: 0.1909830
		}, Vertex{
			x: 0.809017
			y: -0.1909830
			z: -0.1909830
		}, Vertex{
			x: 0.1909830
			y: 0.1909830
			z: -0.809017
		}, Vertex{
			x: 0.1909830
			y: 0.1909830
			z: 0.809017
		}, Vertex{
			x: -0.1909830
			y: 0.1909830
			z: -0.809017
		}, Vertex{
			x: -0.1909830
			y: 0.1909830
			z: 0.809017
		}, Vertex{
			x: 0.1909830
			y: -0.1909830
			z: -0.809017
		}, Vertex{
			x: 0.1909830
			y: -0.1909830
			z: 0.809017
		}, Vertex{
			x: -0.1909830
			y: -0.1909830
			z: -0.809017
		}, Vertex{
			x: -0.1909830
			y: -0.1909830
			z: 0.809017
		}, Vertex{
			x: 0.1909830
			y: -0.809017
			z: 0.1909830
		}, Vertex{
			x: 0.1909830
			y: -0.809017
			z: -0.1909830
		}, Vertex{
			x: -0.1909830
			y: -0.809017
			z: 0.1909830
		}, Vertex{
			x: -0.1909830
			y: -0.809017
			z: -0.1909830
		}, Vertex{
			x: 0.1909830
			y: 0.809017
			z: 0.1909830
		}, Vertex{
			x: 0.1909830
			y: 0.809017
			z: -0.1909830
		}, Vertex{
			x: -0.1909830
			y: 0.809017
			z: 0.1909830
		}, Vertex{
			x: -0.1909830
			y: 0.809017
			z: -0.1909830
		}]
		faces:     [[0, 2, 42, 26, 51, 35, 31, 47, 22, 38], [1, 3, 41, 25, 48, 32, 28, 44, 21, 37],
			[2, 0, 36, 20, 45, 29, 33, 49, 24, 40], [3, 1, 39, 23, 46, 30, 34, 50, 27, 43],
			[4, 5, 47, 31, 59, 19, 17, 57, 29, 45], [5, 4, 44, 28, 56, 16, 18, 58, 30, 46],
			[6, 7, 50, 34, 54, 14, 12, 52, 32, 48], [7, 6, 49, 33, 53, 13, 15, 55, 35, 51],
			[8, 9, 57, 17, 43, 27, 26, 42, 16, 56], [9, 8, 52, 12, 38, 22, 23, 39, 13, 53],
			[10, 11, 55, 15, 37, 21, 20, 36, 14, 54], [11, 10, 58, 18, 40, 24, 25, 41, 19, 59],
			[0, 38, 12, 14, 36], [1, 37, 15, 13, 39], [2, 40, 18, 16, 42],
			[3, 43, 17, 19, 41], [4, 45, 20, 21, 44], [5, 46, 23, 22, 47],
			[6, 48, 25, 24, 49], [7, 51, 26, 27, 50], [8, 56, 28, 32, 52],
			[9, 53, 33, 29, 57], [10, 54, 34, 30, 58], [11, 59, 31, 35, 55]]
	},
	Polyhedron{
		name:      'TruncatedDodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.309017
			y: 0.1909830
			z: 1.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: -1.618034
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: 1.618034
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: -1.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: 1.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: -1.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: 1.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: -1.618034
		}, Vertex{
			x: 1.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: 1.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: 1.618034
			y: -0.309017
			z: 0.1909830
		}, Vertex{
			x: 1.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: -1.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: -1.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: -1.618034
			y: -0.309017
			z: 0.1909830
		}, Vertex{
			x: -1.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.1909830
			y: 1.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: 1.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: -1.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: -1.618034
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: 1.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: 1.618034
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: -1.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: -1.618034
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 1.5
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.5
		}, Vertex{
			x: 1.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.5
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.5
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.5
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 1.0
			z: 1.309017
		}, Vertex{
			x: 0.1909830
			y: 1.0
			z: -1.309017
		}, Vertex{
			x: 0.1909830
			y: -1.0
			z: 1.309017
		}, Vertex{
			x: 0.1909830
			y: -1.0
			z: -1.309017
		}, Vertex{
			x: -0.1909830
			y: 1.0
			z: 1.309017
		}, Vertex{
			x: -0.1909830
			y: 1.0
			z: -1.309017
		}, Vertex{
			x: -0.1909830
			y: -1.0
			z: 1.309017
		}, Vertex{
			x: -0.1909830
			y: -1.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.1909830
			z: 1.0
		}, Vertex{
			x: 1.309017
			y: 0.1909830
			z: -1.0
		}, Vertex{
			x: 1.309017
			y: -0.1909830
			z: 1.0
		}, Vertex{
			x: 1.309017
			y: -0.1909830
			z: -1.0
		}, Vertex{
			x: -1.309017
			y: 0.1909830
			z: 1.0
		}, Vertex{
			x: -1.309017
			y: 0.1909830
			z: -1.0
		}, Vertex{
			x: -1.309017
			y: -0.1909830
			z: 1.0
		}, Vertex{
			x: -1.309017
			y: -0.1909830
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 1.309017
			z: 0.1909830
		}, Vertex{
			x: 1.0
			y: 1.309017
			z: -0.1909830
		}, Vertex{
			x: 1.0
			y: -1.309017
			z: 0.1909830
		}, Vertex{
			x: 1.0
			y: -1.309017
			z: -0.1909830
		}, Vertex{
			x: -1.0
			y: 1.309017
			z: 0.1909830
		}, Vertex{
			x: -1.0
			y: 1.309017
			z: -0.1909830
		}, Vertex{
			x: -1.0
			y: -1.309017
			z: 0.1909830
		}, Vertex{
			x: -1.0
			y: -1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.809017
			y: 0.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: 0.618034
			z: -1.309017
		}, Vertex{
			x: 0.809017
			y: -0.618034
			z: 1.309017
		}, Vertex{
			x: 0.809017
			y: -0.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: 0.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: 0.618034
			z: -1.309017
		}, Vertex{
			x: -0.809017
			y: -0.618034
			z: 1.309017
		}, Vertex{
			x: -0.809017
			y: -0.618034
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: 0.618034
		}, Vertex{
			x: 1.309017
			y: 0.809017
			z: -0.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: 0.618034
		}, Vertex{
			x: 1.309017
			y: -0.809017
			z: -0.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: 0.618034
		}, Vertex{
			x: -1.309017
			y: 0.809017
			z: -0.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: 0.618034
		}, Vertex{
			x: -1.309017
			y: -0.809017
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: 0.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: 0.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: 0.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: -0.618034
			y: 1.309017
			z: 0.809017
		}, Vertex{
			x: -0.618034
			y: 1.309017
			z: -0.809017
		}, Vertex{
			x: -0.618034
			y: -1.309017
			z: 0.809017
		}, Vertex{
			x: -0.618034
			y: -1.309017
			z: -0.809017
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: -0.5
		}]
		faces:     [[0, 74, 56, 24, 26, 58, 72, 2, 106, 104],
			[1, 105, 107, 3, 73, 59, 27, 25, 57, 75], [4, 108, 110, 6, 76, 62, 30, 28, 60, 78],
			[5, 79, 61, 29, 31, 63, 77, 7, 111, 109], [8, 81, 64, 32, 33, 65, 80, 9, 113, 112],
			[10, 114, 115, 11, 82, 67, 35, 34, 66, 83], [12, 116, 117, 13, 84, 69, 37, 36, 68, 85],
			[14, 87, 70, 38, 39, 71, 86, 15, 119, 118], [16, 92, 48, 40, 44, 52, 88, 20, 100, 96],
			[17, 97, 101, 21, 89, 53, 45, 41, 49, 93], [18, 98, 102, 22, 90, 54, 46, 42, 50, 94],
			[19, 95, 51, 43, 47, 55, 91, 23, 103, 99], [0, 52, 44, 45, 53, 1, 75, 115, 114, 74],
			[2, 72, 112, 113, 73, 3, 55, 47, 46, 54], [4, 78, 118, 119, 79, 5, 49, 41, 40, 48],
			[6, 50, 42, 43, 51, 7, 77, 117, 116, 76], [8, 58, 26, 30, 62, 12, 85, 101, 97, 81],
			[9, 80, 96, 100, 84, 13, 63, 31, 27, 59], [10, 83, 99, 103, 87, 14, 60, 28, 24, 56],
			[11, 57, 25, 29, 61, 15, 86, 102, 98, 82], [16, 65, 33, 35, 67, 18, 94, 110, 108, 92],
			[17, 93, 109, 111, 95, 19, 66, 34, 32, 64], [20, 88, 104, 106, 90, 22, 71, 39, 37, 69],
			[21, 68, 36, 38, 70, 23, 91, 107, 105, 89], [0, 104, 88, 52],
			[1, 53, 89, 105], [2, 54, 90, 106], [3, 107, 91, 55],
			[4, 48, 92, 108], [5, 109, 93, 49], [6, 110, 94, 50],
			[7, 51, 95, 111], [8, 112, 72, 58], [9, 59, 73, 113],
			[10, 56, 74, 114], [11, 115, 75, 57], [12, 62, 76, 116],
			[13, 117, 77, 63], [14, 118, 78, 60], [15, 61, 79, 119],
			[16, 96, 80, 65], [17, 64, 81, 97], [18, 67, 82, 98],
			[19, 99, 83, 66], [20, 69, 84, 100], [21, 101, 85, 68],
			[22, 102, 86, 71], [23, 70, 87, 103], [24, 28, 30, 26],
			[25, 27, 31, 29], [32, 34, 35, 33], [36, 37, 39, 38],
			[40, 41, 45, 44], [42, 46, 47, 43]]
	},
	Polyhedron{
		name:      'Icosidodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.1909830
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: 1.0
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: -1.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: 1.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: -1.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: 1.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: -1.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: 1.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: 1.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: 1.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: 1.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: -1.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: -1.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: -1.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: -1.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: 1.0
			z: -0.309017
		}, Vertex{
			x: 0.809017
			y: -1.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: -1.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: 1.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: 1.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: -1.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: -1.0
			z: -0.309017
		}]
		faces:     [[0, 42, 10, 55, 5, 44], [0, 46, 4, 53, 8, 40],
			[2, 36, 8, 57, 6, 50], [2, 48, 7, 59, 10, 38], [15, 13, 53, 20, 22, 55],
			[15, 19, 49, 33, 29, 45], [17, 13, 47, 31, 35, 51],
			[17, 19, 59, 26, 24, 57], [30, 46, 12, 16, 50, 34],
			[30, 42, 26, 27, 43, 31], [32, 48, 18, 14, 44, 28],
			[32, 36, 20, 21, 37, 33], [39, 23, 22, 38, 34, 35],
			[39, 11, 58, 7, 49, 3], [41, 25, 24, 40, 28, 29],
			[41, 9, 52, 4, 47, 1], [54, 11, 43, 1, 45, 5], [54, 23, 21, 52, 12, 14],
			[56, 9, 37, 3, 51, 6], [56, 25, 27, 58, 18, 16], [0, 40, 24, 26, 42],
			[1, 43, 27, 25, 41], [2, 38, 22, 20, 36], [3, 37, 21, 23, 39],
			[4, 46, 30, 31, 47], [5, 45, 29, 28, 44], [6, 51, 35, 34, 50],
			[7, 48, 32, 33, 49], [8, 53, 13, 17, 57], [9, 56, 16, 12, 52],
			[10, 59, 19, 15, 55], [11, 54, 14, 18, 58], [0, 44, 14, 12, 46],
			[1, 47, 13, 15, 45], [2, 50, 16, 18, 48], [3, 49, 19, 17, 51],
			[4, 52, 21, 20, 53], [5, 55, 22, 23, 54], [6, 57, 24, 25, 56],
			[7, 58, 27, 26, 59], [8, 36, 32, 28, 40], [9, 41, 29, 33, 37],
			[10, 42, 30, 34, 38], [11, 39, 35, 31, 43]]
	},
	Polyhedron{
		name:      'GreatDodecicosidodecahedron'
		vertexes_: [Vertex{
			x: -0.5
			y: -0.5
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: 0.1909830
		}, Vertex{
			x: -0.690983
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.309017
			y: -0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: 0.618034
		}, Vertex{
			x: -0.309017
			y: -0.1909830
			z: -0.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: 0.618034
		}, Vertex{
			x: 0.309017
			y: 0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: 0.618034
		}, Vertex{
			x: -0.309017
			y: 0.1909830
			z: -0.618034
		}, Vertex{
			x: -0.1909830
			y: 0.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: 0.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: 0.618034
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: -0.618034
			z: 0.309017
		}, Vertex{
			x: -0.1909830
			y: -0.618034
			z: -0.309017
		}, Vertex{
			x: 0.1909830
			y: -0.618034
			z: 0.309017
		}, Vertex{
			x: 0.1909830
			y: -0.618034
			z: -0.309017
		}, Vertex{
			x: 0.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: -0.618034
			y: 0.309017
			z: -0.1909830
		}, Vertex{
			x: -0.618034
			y: 0.309017
			z: 0.1909830
		}, Vertex{
			x: 0.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: 0.618034
			y: -0.309017
			z: 0.1909830
		}, Vertex{
			x: -0.618034
			y: -0.309017
			z: -0.1909830
		}, Vertex{
			x: -0.618034
			y: -0.309017
			z: 0.1909830
		}]
		faces:     [[0, 24, 56, 48, 12, 14, 50, 58, 26, 2], [0, 36, 44, 32, 17, 21, 34, 48, 40,
			4],
			[7, 3, 39, 47, 33, 18, 22, 35, 51, 43], [7, 5, 25, 53, 45, 9, 11, 47, 55, 27],
			[10, 8, 44, 52, 24, 4, 6, 26, 54, 46], [10, 11, 29, 37, 53, 17, 16, 52, 36, 28],
			[13, 31, 43, 59, 23, 22, 58, 42, 30, 12], [13, 49, 57, 25, 1, 3, 27, 59, 51, 15],
			[19, 33, 46, 38, 2, 6, 42, 50, 35, 23], [19, 55, 39, 29, 9, 8, 28, 38, 54, 18],
			[20, 16, 32, 45, 37, 1, 5, 41, 49, 34], [20, 21, 57, 41, 31, 15, 14, 30, 40, 56],
			[24, 52, 16, 20, 56], [25, 57, 21, 17, 53], [26, 58, 22, 18, 54],
			[27, 55, 19, 23, 59], [28, 36, 0, 2, 38], [29, 39, 3, 1, 37],
			[30, 42, 6, 4, 40], [31, 41, 5, 7, 43], [32, 44, 8, 9, 45],
			[33, 47, 11, 10, 46], [34, 49, 13, 12, 48], [35, 50, 14, 15, 51],
			[24, 0, 4], [25, 5, 1], [26, 6, 2], [27, 3, 7], [28, 8, 10],
			[29, 11, 9], [30, 14, 12], [31, 13, 15], [32, 16, 17],
			[33, 19, 18], [34, 21, 20], [35, 22, 23], [36, 52, 44],
			[37, 45, 53], [38, 46, 54], [39, 55, 47], [40, 48, 56],
			[41, 57, 49], [42, 58, 50], [43, 51, 59]]
	},
	Polyhedron{
		name:      'GreatTruncatedIcosidodecahedron'
		vertexes_: [Vertex{
			x: 0.5
			y: 0.5
			z: -0.7360680
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.7360680
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.7360680
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.7360680
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.7360680
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.7360680
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.7360680
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 0.7360680
		}, Vertex{
			x: 0.5
			y: -0.7360680
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.7360680
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.7360680
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.7360680
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.7360680
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.7360680
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.7360680
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.7360680
			z: -0.5
		}, Vertex{
			x: -0.7360680
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.7360680
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.7360680
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 0.7360680
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.7360680
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.7360680
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.7360680
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.7360680
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 1.0
			z: 0.07294902
		}, Vertex{
			x: 0.1909830
			y: 1.0
			z: -0.07294902
		}, Vertex{
			x: -0.1909830
			y: 1.0
			z: 0.07294902
		}, Vertex{
			x: -0.1909830
			y: 1.0
			z: -0.07294902
		}, Vertex{
			x: 0.1909830
			y: -1.0
			z: 0.07294902
		}, Vertex{
			x: 0.1909830
			y: -1.0
			z: -0.07294902
		}, Vertex{
			x: -0.1909830
			y: -1.0
			z: 0.07294902
		}, Vertex{
			x: -0.1909830
			y: -1.0
			z: -0.07294902
		}, Vertex{
			x: 1.0
			y: 0.07294902
			z: 0.1909830
		}, Vertex{
			x: 1.0
			y: 0.07294902
			z: -0.1909830
		}, Vertex{
			x: -1.0
			y: 0.07294902
			z: 0.1909830
		}, Vertex{
			x: -1.0
			y: 0.07294902
			z: -0.1909830
		}, Vertex{
			x: 1.0
			y: -0.07294902
			z: 0.1909830
		}, Vertex{
			x: 1.0
			y: -0.07294902
			z: -0.1909830
		}, Vertex{
			x: -1.0
			y: -0.07294902
			z: 0.1909830
		}, Vertex{
			x: -1.0
			y: -0.07294902
			z: -0.1909830
		}, Vertex{
			x: 0.07294902
			y: 0.1909830
			z: 1.0
		}, Vertex{
			x: 0.07294902
			y: 0.1909830
			z: -1.0
		}, Vertex{
			x: -0.07294902
			y: 0.1909830
			z: 1.0
		}, Vertex{
			x: -0.07294902
			y: 0.1909830
			z: -1.0
		}, Vertex{
			x: 0.07294902
			y: -0.1909830
			z: 1.0
		}, Vertex{
			x: 0.07294902
			y: -0.1909830
			z: -1.0
		}, Vertex{
			x: -0.07294902
			y: -0.1909830
			z: 1.0
		}, Vertex{
			x: -0.07294902
			y: -0.1909830
			z: -1.0
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: 0.881966
		}, Vertex{
			x: -0.1180340
			y: 0.5
			z: -0.881966
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: 0.881966
		}, Vertex{
			x: 0.1180340
			y: 0.5
			z: -0.881966
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: 0.881966
		}, Vertex{
			x: -0.1180340
			y: -0.5
			z: -0.881966
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: 0.881966
		}, Vertex{
			x: 0.1180340
			y: -0.5
			z: -0.881966
		}, Vertex{
			x: 0.5
			y: 0.881966
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: 0.881966
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: 0.881966
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: 0.881966
			z: 0.1180340
		}, Vertex{
			x: 0.5
			y: -0.881966
			z: -0.1180340
		}, Vertex{
			x: 0.5
			y: -0.881966
			z: 0.1180340
		}, Vertex{
			x: -0.5
			y: -0.881966
			z: -0.1180340
		}, Vertex{
			x: -0.5
			y: -0.881966
			z: 0.1180340
		}, Vertex{
			x: 0.881966
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: 0.881966
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: -0.881966
			y: -0.1180340
			z: 0.5
		}, Vertex{
			x: -0.881966
			y: -0.1180340
			z: -0.5
		}, Vertex{
			x: 0.881966
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: 0.881966
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: -0.881966
			y: 0.1180340
			z: 0.5
		}, Vertex{
			x: -0.881966
			y: 0.1180340
			z: -0.5
		}, Vertex{
			x: -0.618034
			y: 0.690983
			z: -0.4270510
		}, Vertex{
			x: -0.618034
			y: 0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.618034
			y: 0.690983
			z: -0.4270510
		}, Vertex{
			x: 0.618034
			y: 0.690983
			z: 0.4270510
		}, Vertex{
			x: -0.618034
			y: -0.690983
			z: -0.4270510
		}, Vertex{
			x: -0.618034
			y: -0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.618034
			y: -0.690983
			z: -0.4270510
		}, Vertex{
			x: 0.618034
			y: -0.690983
			z: 0.4270510
		}, Vertex{
			x: 0.690983
			y: -0.4270510
			z: -0.618034
		}, Vertex{
			x: 0.690983
			y: -0.4270510
			z: 0.618034
		}, Vertex{
			x: -0.690983
			y: -0.4270510
			z: -0.618034
		}, Vertex{
			x: -0.690983
			y: -0.4270510
			z: 0.618034
		}, Vertex{
			x: 0.690983
			y: 0.4270510
			z: -0.618034
		}, Vertex{
			x: 0.690983
			y: 0.4270510
			z: 0.618034
		}, Vertex{
			x: -0.690983
			y: 0.4270510
			z: -0.618034
		}, Vertex{
			x: -0.690983
			y: 0.4270510
			z: 0.618034
		}, Vertex{
			x: -0.4270510
			y: -0.618034
			z: 0.690983
		}, Vertex{
			x: -0.4270510
			y: -0.618034
			z: -0.690983
		}, Vertex{
			x: 0.4270510
			y: -0.618034
			z: 0.690983
		}, Vertex{
			x: 0.4270510
			y: -0.618034
			z: -0.690983
		}, Vertex{
			x: -0.4270510
			y: 0.618034
			z: 0.690983
		}, Vertex{
			x: -0.4270510
			y: 0.618034
			z: -0.690983
		}, Vertex{
			x: 0.4270510
			y: 0.618034
			z: 0.690983
		}, Vertex{
			x: 0.4270510
			y: 0.618034
			z: -0.690983
		}, Vertex{
			x: -0.927051
			y: 0.1909830
			z: 0.3819660
		}, Vertex{
			x: -0.927051
			y: 0.1909830
			z: -0.3819660
		}, Vertex{
			x: 0.927051
			y: 0.1909830
			z: 0.3819660
		}, Vertex{
			x: 0.927051
			y: 0.1909830
			z: -0.3819660
		}, Vertex{
			x: -0.927051
			y: -0.1909830
			z: 0.3819660
		}, Vertex{
			x: -0.927051
			y: -0.1909830
			z: -0.3819660
		}, Vertex{
			x: 0.927051
			y: -0.1909830
			z: 0.3819660
		}, Vertex{
			x: 0.927051
			y: -0.1909830
			z: -0.3819660
		}, Vertex{
			x: 0.1909830
			y: 0.3819660
			z: -0.927051
		}, Vertex{
			x: 0.1909830
			y: 0.3819660
			z: 0.927051
		}, Vertex{
			x: -0.1909830
			y: 0.3819660
			z: -0.927051
		}, Vertex{
			x: -0.1909830
			y: 0.3819660
			z: 0.927051
		}, Vertex{
			x: 0.1909830
			y: -0.3819660
			z: -0.927051
		}, Vertex{
			x: 0.1909830
			y: -0.3819660
			z: 0.927051
		}, Vertex{
			x: -0.1909830
			y: -0.3819660
			z: -0.927051
		}, Vertex{
			x: -0.1909830
			y: -0.3819660
			z: 0.927051
		}, Vertex{
			x: 0.3819660
			y: -0.927051
			z: 0.1909830
		}, Vertex{
			x: 0.3819660
			y: -0.927051
			z: -0.1909830
		}, Vertex{
			x: -0.3819660
			y: -0.927051
			z: 0.1909830
		}, Vertex{
			x: -0.3819660
			y: -0.927051
			z: -0.1909830
		}, Vertex{
			x: 0.3819660
			y: 0.927051
			z: 0.1909830
		}, Vertex{
			x: 0.3819660
			y: 0.927051
			z: -0.1909830
		}, Vertex{
			x: -0.3819660
			y: 0.927051
			z: 0.1909830
		}, Vertex{
			x: -0.3819660
			y: 0.927051
			z: -0.1909830
		}]
		faces:     [[0, 2, 26, 74, 106, 58, 56, 104, 72, 24],
			[1, 25, 73, 105, 57, 59, 107, 75, 27, 3], [4, 28, 76, 108, 60, 62, 110, 78, 30, 6],
			[5, 7, 31, 79, 111, 63, 61, 109, 77, 29], [8, 9, 33, 81, 113, 65, 64, 112, 80, 32],
			[10, 34, 82, 114, 66, 67, 115, 83, 35, 11], [12, 36, 84, 116, 68, 69, 117, 85, 37, 13],
			[14, 15, 39, 87, 119, 71, 70, 118, 86, 38], [16, 20, 44, 92, 100, 52, 48, 96, 88, 40],
			[17, 41, 89, 97, 49, 53, 101, 93, 45, 21], [18, 42, 90, 98, 50, 54, 102, 94, 46, 22],
			[19, 23, 47, 95, 103, 55, 51, 99, 91, 43], [0, 24, 48, 52, 28, 4],
			[1, 5, 29, 53, 49, 25], [2, 6, 30, 54, 50, 26], [3, 27, 51, 55, 31, 7],
			[8, 32, 56, 58, 34, 10], [9, 11, 35, 59, 57, 33],
			[12, 14, 38, 62, 60, 36], [13, 37, 61, 63, 39, 15],
			[16, 40, 64, 65, 41, 17], [18, 19, 43, 67, 66, 42],
			[20, 21, 45, 69, 68, 44], [22, 46, 70, 71, 47, 23],
			[72, 104, 80, 112, 88, 96], [73, 97, 89, 113, 81, 105],
			[74, 98, 90, 114, 82, 106], [75, 107, 83, 115, 91, 99],
			[76, 100, 92, 116, 84, 108], [77, 109, 85, 117, 93, 101],
			[78, 110, 86, 118, 94, 102], [79, 103, 95, 119, 87, 111],
			[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9], [12, 13, 15, 14],
			[16, 17, 21, 20], [18, 22, 23, 19], [24, 72, 96, 48],
			[25, 49, 97, 73], [26, 50, 98, 74], [27, 75, 99, 51],
			[28, 52, 100, 76], [29, 77, 101, 53], [30, 78, 102, 54],
			[31, 55, 103, 79], [32, 80, 104, 56], [33, 57, 105, 81],
			[34, 58, 106, 82], [35, 83, 107, 59], [36, 60, 108, 84],
			[37, 85, 109, 61], [38, 86, 110, 62], [39, 63, 111, 87],
			[40, 88, 112, 64], [41, 65, 113, 89], [42, 66, 114, 90],
			[43, 91, 115, 67], [44, 68, 116, 92], [45, 93, 117, 69],
			[46, 94, 118, 70], [47, 71, 119, 95]]
	},
	Polyhedron{
		name:      'GreatInvertedSnubIcosidodecahedron'
		vertexes_: [Vertex{
			x: -0.4635223
			y: 0.1874755
			z: -0.4074937
		}, Vertex{
			x: 0.4635223
			y: 0.1874755
			z: 0.4074937
		}, Vertex{
			x: 0.4635223
			y: -0.1874755
			z: -0.4074937
		}, Vertex{
			x: -0.4635223
			y: -0.1874755
			z: 0.4074937
		}, Vertex{
			x: -0.1874755
			y: -0.4074937
			z: 0.4635223
		}, Vertex{
			x: 0.1874755
			y: -0.4074937
			z: -0.4635223
		}, Vertex{
			x: 0.1874755
			y: 0.4074937
			z: 0.4635223
		}, Vertex{
			x: -0.1874755
			y: 0.4074937
			z: -0.4635223
		}, Vertex{
			x: 0.4074937
			y: 0.4635223
			z: 0.1874755
		}, Vertex{
			x: -0.4074937
			y: 0.4635223
			z: -0.1874755
		}, Vertex{
			x: -0.4074937
			y: -0.4635223
			z: 0.1874755
		}, Vertex{
			x: 0.4074937
			y: -0.4635223
			z: -0.1874755
		}, Vertex{
			x: 0.2291837
			y: 0.5666434
			z: 0.2060127
		}, Vertex{
			x: -0.2291837
			y: 0.5666434
			z: -0.2060127
		}, Vertex{
			x: -0.2291837
			y: -0.5666434
			z: 0.2060127
		}, Vertex{
			x: 0.2291837
			y: -0.5666434
			z: -0.2060127
		}, Vertex{
			x: 0.5666434
			y: 0.2060127
			z: 0.2291837
		}, Vertex{
			x: -0.5666434
			y: 0.2060127
			z: -0.2291837
		}, Vertex{
			x: -0.5666434
			y: -0.2060127
			z: 0.2291837
		}, Vertex{
			x: 0.5666434
			y: -0.2060127
			z: -0.2291837
		}, Vertex{
			x: 0.2060127
			y: 0.2291837
			z: 0.5666434
		}, Vertex{
			x: -0.2060127
			y: 0.2291837
			z: -0.5666434
		}, Vertex{
			x: -0.2060127
			y: -0.2291837
			z: 0.5666434
		}, Vertex{
			x: 0.2060127
			y: -0.2291837
			z: -0.5666434
		}, Vertex{
			x: -0.1133175
			y: 0.3791678
			z: 0.5093545
		}, Vertex{
			x: 0.1133175
			y: 0.3791678
			z: -0.5093545
		}, Vertex{
			x: 0.1133175
			y: -0.3791678
			z: 0.5093545
		}, Vertex{
			x: -0.1133175
			y: -0.3791678
			z: -0.5093545
		}, Vertex{
			x: -0.3791678
			y: 0.5093545
			z: 0.1133175
		}, Vertex{
			x: 0.3791678
			y: 0.5093545
			z: -0.1133175
		}, Vertex{
			x: 0.3791678
			y: -0.5093545
			z: 0.1133175
		}, Vertex{
			x: -0.3791678
			y: -0.5093545
			z: -0.1133175
		}, Vertex{
			x: -0.5093545
			y: 0.1133175
			z: 0.3791678
		}, Vertex{
			x: 0.5093545
			y: 0.1133175
			z: -0.3791678
		}, Vertex{
			x: 0.5093545
			y: -0.1133175
			z: 0.3791678
		}, Vertex{
			x: -0.5093545
			y: -0.1133175
			z: -0.3791678
		}, Vertex{
			x: 0.5208111
			y: 0.2801708
			z: -0.2575096
		}, Vertex{
			x: -0.5208111
			y: 0.2801708
			z: 0.2575096
		}, Vertex{
			x: -0.5208111
			y: -0.2801708
			z: -0.2575096
		}, Vertex{
			x: 0.5208111
			y: -0.2801708
			z: 0.2575096
		}, Vertex{
			x: -0.2801708
			y: -0.2575096
			z: -0.5208111
		}, Vertex{
			x: 0.2801708
			y: -0.2575096
			z: 0.5208111
		}, Vertex{
			x: 0.2801708
			y: 0.2575096
			z: -0.5208111
		}, Vertex{
			x: -0.2801708
			y: 0.2575096
			z: 0.5208111
		}, Vertex{
			x: 0.2575096
			y: -0.5208111
			z: 0.2801708
		}, Vertex{
			x: -0.2575096
			y: -0.5208111
			z: -0.2801708
		}, Vertex{
			x: -0.2575096
			y: 0.5208111
			z: 0.2801708
		}, Vertex{
			x: 0.2575096
			y: 0.5208111
			z: -0.2801708
		}, Vertex{
			x: 0.09269529
			y: 0.04583221
			z: -0.6366774
		}, Vertex{
			x: -0.09269529
			y: 0.04583221
			z: 0.6366774
		}, Vertex{
			x: -0.09269529
			y: -0.04583221
			z: -0.6366774
		}, Vertex{
			x: 0.09269529
			y: -0.04583221
			z: 0.6366774
		}, Vertex{
			x: 0.04583221
			y: -0.6366774
			z: 0.09269529
		}, Vertex{
			x: -0.04583221
			y: -0.6366774
			z: -0.09269529
		}, Vertex{
			x: -0.04583221
			y: 0.6366774
			z: 0.09269529
		}, Vertex{
			x: 0.04583221
			y: 0.6366774
			z: -0.09269529
		}, Vertex{
			x: -0.6366774
			y: 0.09269529
			z: 0.04583221
		}, Vertex{
			x: 0.6366774
			y: 0.09269529
			z: -0.04583221
		}, Vertex{
			x: 0.6366774
			y: -0.09269529
			z: 0.04583221
		}, Vertex{
			x: -0.6366774
			y: -0.09269529
			z: -0.04583221
		}]
		faces:     [[0, 36, 28, 48, 12], [1, 37, 29, 49, 13],
			[2, 38, 30, 50, 14], [3, 39, 31, 51, 15], [4, 40, 32, 53, 17],
			[5, 41, 33, 52, 16], [6, 42, 34, 55, 19], [7, 43, 35, 54, 18],
			[8, 44, 24, 58, 22], [9, 45, 25, 59, 23], [10, 46, 26, 56, 20],
			[11, 47, 27, 57, 21], [0, 2, 14], [1, 3, 15], [2, 0, 12],
			[3, 1, 13], [4, 5, 16], [5, 4, 17], [6, 7, 18], [7, 6, 19],
			[8, 11, 21], [9, 10, 20], [10, 9, 23], [11, 8, 22],
			[12, 48, 56], [13, 49, 57], [14, 50, 58], [15, 51, 59],
			[16, 52, 48], [17, 53, 49], [18, 54, 50], [19, 55, 51],
			[20, 56, 52], [21, 57, 53], [22, 58, 54], [23, 59, 55],
			[24, 44, 36], [25, 45, 37], [26, 46, 38], [27, 47, 39],
			[28, 36, 40], [29, 37, 41], [30, 38, 42], [31, 39, 43],
			[32, 40, 44], [33, 41, 45], [34, 42, 46], [35, 43, 47],
			[36, 0, 24], [37, 1, 25], [38, 2, 26], [39, 3, 27],
			[40, 4, 28], [41, 5, 29], [42, 6, 30], [43, 7, 31],
			[44, 8, 32], [45, 9, 33], [46, 10, 34], [47, 11, 35],
			[48, 28, 16], [49, 29, 17], [50, 30, 18], [51, 31, 19],
			[52, 33, 20], [53, 32, 21], [54, 35, 22], [55, 34, 23],
			[56, 26, 12], [57, 27, 13], [58, 24, 14], [59, 25, 15],
			[24, 0, 14], [25, 1, 15], [26, 2, 12], [27, 3, 13],
			[28, 4, 16], [29, 5, 17], [30, 6, 18], [31, 7, 19],
			[32, 8, 21], [33, 9, 20], [34, 10, 23], [35, 11, 22],
			[36, 44, 40], [37, 45, 41], [38, 46, 42], [39, 47, 43],
			[48, 52, 56], [49, 53, 57], [50, 54, 58], [51, 55, 59]]
	},
	Polyhedron{
		name:      'DitrigonalDodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: 0.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: 0.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: 0.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: 0.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: 0.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: 0.0
			z: -0.309017
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: 0.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.5
		}]
		faces:     [[0, 6, 2, 16, 18], [0, 8, 16, 12, 10], [0, 14, 12, 2, 4],
			[7, 1, 19, 17, 3], [7, 11, 6, 19, 18], [7, 16, 17, 6, 10],
			[9, 2, 11, 14, 18], [9, 5, 14, 15, 4], [9, 19, 15, 11, 3],
			[13, 12, 5, 8, 4], [13, 15, 1, 5, 3], [13, 17, 8, 1, 10],
			[0, 4, 15, 19, 6], [0, 10, 1, 15, 14], [0, 18, 19, 1, 8],
			[7, 3, 5, 12, 16], [7, 10, 12, 14, 11], [7, 18, 14, 5, 1],
			[9, 3, 17, 16, 2], [9, 4, 8, 17, 19], [9, 18, 16, 8, 5],
			[13, 3, 11, 2, 12], [13, 4, 2, 6, 17], [13, 10, 6, 11, 15]]
	},
	Polyhedron{
		name:      'MedialDisdyakisTriacontahedron'
		vertexes_: [Vertex{
			x: 3.618034
			y: 0.0
			z: 5.854102
		}, Vertex{
			x: 3.618034
			y: 0.0
			z: -5.854102
		}, Vertex{
			x: -3.618034
			y: 0.0
			z: 5.854102
		}, Vertex{
			x: -3.618034
			y: 0.0
			z: -5.854102
		}, Vertex{
			x: 5.854102
			y: 3.618034
			z: 0.0
		}, Vertex{
			x: 5.854102
			y: -3.618034
			z: 0.0
		}, Vertex{
			x: -5.854102
			y: 3.618034
			z: 0.0
		}, Vertex{
			x: -5.854102
			y: -3.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 5.854102
			z: 3.618034
		}, Vertex{
			x: 0.0
			y: 5.854102
			z: -3.618034
		}, Vertex{
			x: 0.0
			y: -5.854102
			z: 3.618034
		}, Vertex{
			x: 0.0
			y: -5.854102
			z: -3.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.666667
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.666667
		}, Vertex{
			x: 1.666667
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.666667
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.666667
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.666667
			z: 0.0
		}, Vertex{
			x: 0.8541020
			y: 0.0
			z: 1.381966
		}, Vertex{
			x: 0.8541020
			y: 0.0
			z: -1.381966
		}, Vertex{
			x: -0.8541020
			y: 0.0
			z: 1.381966
		}, Vertex{
			x: -0.8541020
			y: 0.0
			z: -1.381966
		}, Vertex{
			x: 1.381966
			y: 0.8541020
			z: 0.0
		}, Vertex{
			x: 1.381966
			y: -0.8541020
			z: 0.0
		}, Vertex{
			x: -1.381966
			y: 0.8541020
			z: 0.0
		}, Vertex{
			x: -1.381966
			y: -0.8541020
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.381966
			z: 0.8541020
		}, Vertex{
			x: 0.0
			y: 1.381966
			z: -0.8541020
		}, Vertex{
			x: 0.0
			y: -1.381966
			z: 0.8541020
		}, Vertex{
			x: 0.0
			y: -1.381966
			z: -0.8541020
		}, Vertex{
			x: 0.5150283
			y: 0.8333333
			z: 1.348362
		}, Vertex{
			x: 0.5150283
			y: 0.8333333
			z: -1.348362
		}, Vertex{
			x: 0.5150283
			y: -0.8333333
			z: 1.348362
		}, Vertex{
			x: 0.5150283
			y: -0.8333333
			z: -1.348362
		}, Vertex{
			x: -0.5150283
			y: 0.8333333
			z: 1.348362
		}, Vertex{
			x: -0.5150283
			y: 0.8333333
			z: -1.348362
		}, Vertex{
			x: -0.5150283
			y: -0.8333333
			z: 1.348362
		}, Vertex{
			x: -0.5150283
			y: -0.8333333
			z: -1.348362
		}, Vertex{
			x: 1.348362
			y: 0.5150283
			z: 0.8333333
		}, Vertex{
			x: 1.348362
			y: 0.5150283
			z: -0.8333333
		}, Vertex{
			x: 1.348362
			y: -0.5150283
			z: 0.8333333
		}, Vertex{
			x: 1.348362
			y: -0.5150283
			z: -0.8333333
		}, Vertex{
			x: -1.348362
			y: 0.5150283
			z: 0.8333333
		}, Vertex{
			x: -1.348362
			y: 0.5150283
			z: -0.8333333
		}, Vertex{
			x: -1.348362
			y: -0.5150283
			z: 0.8333333
		}, Vertex{
			x: -1.348362
			y: -0.5150283
			z: -0.8333333
		}, Vertex{
			x: 0.8333333
			y: 1.348362
			z: 0.5150283
		}, Vertex{
			x: 0.8333333
			y: 1.348362
			z: -0.5150283
		}, Vertex{
			x: 0.8333333
			y: -1.348362
			z: 0.5150283
		}, Vertex{
			x: 0.8333333
			y: -1.348362
			z: -0.5150283
		}, Vertex{
			x: -0.8333333
			y: 1.348362
			z: 0.5150283
		}, Vertex{
			x: -0.8333333
			y: 1.348362
			z: -0.5150283
		}, Vertex{
			x: -0.8333333
			y: -1.348362
			z: 0.5150283
		}, Vertex{
			x: -0.8333333
			y: -1.348362
			z: -0.5150283
		}]
		faces:     [[0, 14, 22], [0, 22, 46], [0, 46, 26], [0, 26, 34],
			[0, 34, 20], [0, 20, 36], [0, 36, 28], [0, 28, 48],
			[0, 48, 23], [0, 23, 14], [1, 14, 23], [1, 23, 49],
			[1, 49, 29], [1, 29, 37], [1, 37, 21], [1, 21, 35],
			[1, 35, 27], [1, 27, 47], [1, 47, 22], [1, 22, 14],
			[2, 15, 25], [2, 25, 52], [2, 52, 28], [2, 28, 32],
			[2, 32, 18], [2, 18, 30], [2, 30, 26], [2, 26, 50],
			[2, 50, 24], [2, 24, 15], [3, 15, 24], [3, 24, 51],
			[3, 51, 27], [3, 27, 31], [3, 31, 19], [3, 19, 33],
			[3, 33, 29], [3, 29, 53], [3, 53, 25], [3, 25, 15],
			[4, 16, 26], [4, 26, 30], [4, 30, 18], [4, 18, 40],
			[4, 40, 23], [4, 23, 41], [4, 41, 19], [4, 19, 31],
			[4, 31, 27], [4, 27, 16], [5, 17, 29], [5, 29, 33],
			[5, 33, 19], [5, 19, 39], [5, 39, 22], [5, 22, 38],
			[5, 38, 18], [5, 18, 32], [5, 32, 28], [5, 28, 17],
			[6, 16, 27], [6, 27, 35], [6, 35, 21], [6, 21, 45],
			[6, 45, 25], [6, 25, 44], [6, 44, 20], [6, 20, 34],
			[6, 34, 26], [6, 26, 16], [7, 17, 28], [7, 28, 36],
			[7, 36, 20], [7, 20, 42], [7, 42, 24], [7, 24, 43],
			[7, 43, 21], [7, 21, 37], [7, 37, 29], [7, 29, 17],
			[8, 12, 18], [8, 18, 38], [8, 38, 22], [8, 22, 47],
			[8, 47, 27], [8, 27, 51], [8, 51, 24], [8, 24, 42],
			[8, 42, 20], [8, 20, 12], [9, 13, 21], [9, 21, 43],
			[9, 43, 24], [9, 24, 50], [9, 50, 26], [9, 26, 46],
			[9, 46, 22], [9, 22, 39], [9, 39, 19], [9, 19, 13],
			[10, 12, 20], [10, 20, 44], [10, 44, 25], [10, 25, 53],
			[10, 53, 29], [10, 29, 49], [10, 49, 23], [10, 23, 40],
			[10, 40, 18], [10, 18, 12], [11, 13, 19], [11, 19, 41],
			[11, 41, 23], [11, 23, 48], [11, 48, 28], [11, 28, 52],
			[11, 52, 25], [11, 25, 45], [11, 45, 21], [11, 21, 13]]
	},
	Polyhedron{
		name:      'GreatCubicuboctahedron'
		vertexes_: [Vertex{
			x: -0.5
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -0.2071068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 0.2071068
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -0.2071068
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 0.2071068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -0.2071068
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -0.2071068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.2071068
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -0.2071068
			z: 0.5
		}]
		faces:     [[0, 2, 18, 19, 3, 1, 17, 16], [0, 8, 9, 1, 5, 13, 12, 4],
			[11, 10, 2, 6, 14, 15, 7, 3], [11, 19, 23, 15, 13, 21, 17, 9],
			[20, 12, 14, 22, 18, 10, 8, 16], [20, 21, 5, 7, 23, 22, 6, 4],
			[0, 4, 6, 2], [1, 3, 7, 5], [8, 10, 11, 9], [12, 13, 15, 14],
			[16, 17, 21, 20], [18, 22, 23, 19], [0, 16, 8], [1, 9, 17],
			[2, 10, 18], [3, 19, 11], [4, 12, 20], [5, 21, 13],
			[6, 22, 14], [7, 15, 23]]
	},
	Polyhedron{
		name:      'SmallTriambicIcosahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.2763932
			z: 0.7236068
		}, Vertex{
			x: 0.0
			y: 0.2763932
			z: -0.7236068
		}, Vertex{
			x: 0.0
			y: -0.2763932
			z: 0.7236068
		}, Vertex{
			x: 0.0
			y: -0.2763932
			z: -0.7236068
		}, Vertex{
			x: 0.7236068
			y: 0.0
			z: 0.2763932
		}, Vertex{
			x: 0.7236068
			y: 0.0
			z: -0.2763932
		}, Vertex{
			x: -0.7236068
			y: 0.0
			z: 0.2763932
		}, Vertex{
			x: -0.7236068
			y: 0.0
			z: -0.2763932
		}, Vertex{
			x: 0.2763932
			y: 0.7236068
			z: 0.0
		}, Vertex{
			x: 0.2763932
			y: -0.7236068
			z: 0.0
		}, Vertex{
			x: -0.2763932
			y: 0.7236068
			z: 0.0
		}, Vertex{
			x: -0.2763932
			y: -0.7236068
			z: 0.0
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: -0.3819660
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 0.3819660
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: -0.3819660
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: -0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 0.3819660
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: -0.3819660
		}, Vertex{
			x: 0.4472136
			y: 0.4472136
			z: 0.4472136
		}, Vertex{
			x: 0.4472136
			y: 0.4472136
			z: -0.4472136
		}, Vertex{
			x: 0.4472136
			y: -0.4472136
			z: 0.4472136
		}, Vertex{
			x: 0.4472136
			y: -0.4472136
			z: -0.4472136
		}, Vertex{
			x: -0.4472136
			y: 0.4472136
			z: 0.4472136
		}, Vertex{
			x: -0.4472136
			y: 0.4472136
			z: -0.4472136
		}, Vertex{
			x: -0.4472136
			y: -0.4472136
			z: 0.4472136
		}, Vertex{
			x: -0.4472136
			y: -0.4472136
			z: -0.4472136
		}]
		faces:     [[12, 0, 14, 30, 22, 26], [12, 26, 17, 5, 16, 24],
			[12, 24, 20, 28, 14, 2], [12, 2, 22, 9, 17, 4], [12, 4, 16, 8, 20, 0],
			[15, 1, 13, 27, 23, 31], [15, 31, 19, 6, 18, 29],
			[15, 29, 21, 25, 13, 3], [15, 3, 23, 11, 19, 7], [15, 7, 18, 10, 21, 1],
			[13, 1, 21, 8, 16, 5], [13, 5, 17, 9, 23, 3], [13, 25, 16, 4, 17, 27],
			[14, 0, 20, 10, 18, 6], [14, 6, 19, 11, 22, 2], [14, 28, 18, 7, 19, 30],
			[20, 8, 21, 29, 18, 28], [20, 24, 16, 25, 21, 10],
			[22, 11, 23, 27, 17, 26], [22, 30, 19, 31, 23, 9]]
	},
	Polyhedron{
		name:      'GreatIcosahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: -0.5
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: 0.5
		}]
		faces:     [[0, 2, 10], [0, 10, 5], [0, 5, 4], [0, 4, 8],
			[0, 8, 2], [3, 1, 11], [3, 11, 7], [3, 7, 6], [3, 6, 9],
			[3, 9, 1], [2, 6, 7], [2, 7, 10], [10, 7, 11], [10, 11, 5],
			[5, 11, 1], [5, 1, 4], [4, 1, 9], [4, 9, 8], [8, 9, 6],
			[8, 6, 2]]
	},
	Polyhedron{
		name:      'SmallHexagrammicHexecontahedron'
		vertexes_: [Vertex{
			x: 0.309017
			y: 0.0
			z: -1.366760
		}, Vertex{
			x: 0.309017
			y: 0.0
			z: 1.366760
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: -1.366760
		}, Vertex{
			x: -0.309017
			y: 0.0
			z: 1.366760
		}, Vertex{
			x: -1.366760
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: -1.366760
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: 1.366760
			y: 0.309017
			z: 0.0
		}, Vertex{
			x: 1.366760
			y: -0.309017
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.366760
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: -1.366760
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: 1.366760
			z: 0.309017
		}, Vertex{
			x: 0.0
			y: 1.366760
			z: -0.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: 0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: 1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 0.0
			y: -0.5
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: 0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: -1.309017
			y: 0.0
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: 0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: 1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -0.5
			y: -1.309017
			z: 0.0
		}, Vertex{
			x: -0.2678437
			y: -0.9333802
			z: -1.010241
		}, Vertex{
			x: -0.2678437
			y: -0.9333802
			z: 1.010241
		}, Vertex{
			x: -0.2678437
			y: 0.9333802
			z: -1.010241
		}, Vertex{
			x: -0.2678437
			y: 0.9333802
			z: 1.010241
		}, Vertex{
			x: 0.2678437
			y: -0.9333802
			z: -1.010241
		}, Vertex{
			x: 0.2678437
			y: -0.9333802
			z: 1.010241
		}, Vertex{
			x: 0.2678437
			y: 0.9333802
			z: -1.010241
		}, Vertex{
			x: 0.2678437
			y: 0.9333802
			z: 1.010241
		}, Vertex{
			x: -1.010241
			y: -0.2678437
			z: -0.9333802
		}, Vertex{
			x: -1.010241
			y: -0.2678437
			z: 0.9333802
		}, Vertex{
			x: -1.010241
			y: 0.2678437
			z: -0.9333802
		}, Vertex{
			x: -1.010241
			y: 0.2678437
			z: 0.9333802
		}, Vertex{
			x: 1.010241
			y: -0.2678437
			z: -0.9333802
		}, Vertex{
			x: 1.010241
			y: -0.2678437
			z: 0.9333802
		}, Vertex{
			x: 1.010241
			y: 0.2678437
			z: -0.9333802
		}, Vertex{
			x: 1.010241
			y: 0.2678437
			z: 0.9333802
		}, Vertex{
			x: -0.9333802
			y: -1.010241
			z: -0.2678437
		}, Vertex{
			x: -0.9333802
			y: -1.010241
			z: 0.2678437
		}, Vertex{
			x: -0.9333802
			y: 1.010241
			z: -0.2678437
		}, Vertex{
			x: -0.9333802
			y: 1.010241
			z: 0.2678437
		}, Vertex{
			x: 0.9333802
			y: -1.010241
			z: -0.2678437
		}, Vertex{
			x: 0.9333802
			y: -1.010241
			z: 0.2678437
		}, Vertex{
			x: 0.9333802
			y: 1.010241
			z: -0.2678437
		}, Vertex{
			x: 0.9333802
			y: 1.010241
			z: 0.2678437
		}, Vertex{
			x: -0.1859145
			y: 0.0
			z: -0.3008159
		}, Vertex{
			x: -0.1859145
			y: 0.0
			z: 0.3008159
		}, Vertex{
			x: 0.1859145
			y: 0.0
			z: -0.3008159
		}, Vertex{
			x: 0.1859145
			y: 0.0
			z: 0.3008159
		}, Vertex{
			x: -0.3008159
			y: -0.1859145
			z: 0.0
		}, Vertex{
			x: -0.3008159
			y: 0.1859145
			z: 0.0
		}, Vertex{
			x: 0.3008159
			y: -0.1859145
			z: 0.0
		}, Vertex{
			x: 0.3008159
			y: 0.1859145
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.3008159
			z: -0.1859145
		}, Vertex{
			x: 0.0
			y: -0.3008159
			z: 0.1859145
		}, Vertex{
			x: 0.0
			y: 0.3008159
			z: -0.1859145
		}, Vertex{
			x: 0.0
			y: 0.3008159
			z: 0.1859145
		}, Vertex{
			x: -0.5768607
			y: -0.4333802
			z: -1.201224
		}, Vertex{
			x: -0.5768607
			y: -0.4333802
			z: 1.201224
		}, Vertex{
			x: -0.5768607
			y: 0.4333802
			z: -1.201224
		}, Vertex{
			x: -0.5768607
			y: 0.4333802
			z: 1.201224
		}, Vertex{
			x: 0.5768607
			y: -0.4333802
			z: -1.201224
		}, Vertex{
			x: 0.5768607
			y: -0.4333802
			z: 1.201224
		}, Vertex{
			x: 0.5768607
			y: 0.4333802
			z: -1.201224
		}, Vertex{
			x: 0.5768607
			y: 0.4333802
			z: 1.201224
		}, Vertex{
			x: -1.201224
			y: -0.5768607
			z: -0.4333802
		}, Vertex{
			x: -1.201224
			y: -0.5768607
			z: 0.4333802
		}, Vertex{
			x: -1.201224
			y: 0.5768607
			z: -0.4333802
		}, Vertex{
			x: -1.201224
			y: 0.5768607
			z: 0.4333802
		}, Vertex{
			x: 1.201224
			y: -0.5768607
			z: -0.4333802
		}, Vertex{
			x: 1.201224
			y: -0.5768607
			z: 0.4333802
		}, Vertex{
			x: 1.201224
			y: 0.5768607
			z: -0.4333802
		}, Vertex{
			x: 1.201224
			y: 0.5768607
			z: 0.4333802
		}, Vertex{
			x: -0.4333802
			y: -1.201224
			z: -0.5768607
		}, Vertex{
			x: -0.4333802
			y: -1.201224
			z: 0.5768607
		}, Vertex{
			x: -0.4333802
			y: 1.201224
			z: -0.5768607
		}, Vertex{
			x: -0.4333802
			y: 1.201224
			z: 0.5768607
		}, Vertex{
			x: 0.4333802
			y: -1.201224
			z: -0.5768607
		}, Vertex{
			x: 0.4333802
			y: -1.201224
			z: 0.5768607
		}, Vertex{
			x: 0.4333802
			y: 1.201224
			z: -0.5768607
		}, Vertex{
			x: 0.4333802
			y: 1.201224
			z: 0.5768607
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: 0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: 0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: -0.809017
		}, Vertex{
			x: -0.809017
			y: -0.809017
			z: -0.809017
		}]
		faces:     [[60, 0, 17, 74, 100, 82], [60, 82, 20, 44, 97, 36],
			[60, 36, 12, 2, 16, 38], [60, 38, 101, 46, 21, 80],
			[60, 80, 96, 72, 13, 0], [61, 1, 15, 73, 98, 81],
			[61, 81, 22, 47, 103, 39], [61, 39, 18, 3, 14, 37],
			[61, 37, 99, 45, 23, 83], [61, 83, 102, 75, 19, 1],
			[62, 2, 12, 76, 104, 84], [62, 84, 25, 50, 109, 42],
			[62, 42, 17, 0, 13, 40], [62, 40, 105, 48, 24, 86],
			[62, 86, 108, 78, 16, 2], [63, 3, 18, 79, 110, 87],
			[63, 87, 27, 49, 107, 41], [63, 41, 15, 1, 19, 43],
			[63, 43, 111, 51, 26, 85], [63, 85, 106, 77, 14, 3],
			[64, 4, 22, 81, 98, 89], [64, 89, 29, 52, 97, 44],
			[64, 44, 20, 5, 23, 45], [64, 45, 99, 53, 28, 88],
			[64, 88, 96, 80, 21, 4], [65, 5, 20, 82, 100, 90],
			[65, 90, 31, 55, 103, 47], [65, 47, 22, 4, 21, 46],
			[65, 46, 101, 54, 30, 91], [65, 91, 102, 83, 23, 5],
			[66, 6, 25, 84, 104, 92], [66, 92, 32, 57, 107, 49],
			[66, 49, 27, 7, 24, 48], [66, 48, 105, 56, 33, 93],
			[66, 93, 106, 85, 26, 6], [67, 7, 27, 87, 110, 95],
			[67, 95, 34, 58, 109, 50], [67, 50, 25, 6, 26, 51],
			[67, 51, 111, 59, 35, 94], [67, 94, 108, 86, 24, 7],
			[68, 8, 32, 92, 104, 76], [68, 76, 12, 36, 97, 52],
			[68, 52, 29, 9, 33, 56], [68, 56, 105, 40, 13, 72],
			[68, 72, 96, 88, 28, 8], [69, 9, 29, 89, 98, 73],
			[69, 73, 15, 41, 107, 57], [69, 57, 32, 8, 28, 53],
			[69, 53, 99, 37, 14, 77], [69, 77, 106, 93, 33, 9],
			[70, 10, 31, 90, 100, 74], [70, 74, 17, 42, 109, 58],
			[70, 58, 34, 11, 30, 54], [70, 54, 101, 38, 16, 78],
			[70, 78, 108, 94, 35, 10], [71, 11, 34, 95, 110, 79],
			[71, 79, 18, 39, 103, 55], [71, 55, 31, 10, 35, 59],
			[71, 59, 111, 43, 19, 75], [71, 75, 102, 91, 30, 11]]
	},
	Polyhedron{
		name:      'TridyakisIcosahedron'
		vertexes_: [Vertex{
			x: 1.677051
			y: 0.0
			z: 2.713526
		}, Vertex{
			x: 1.677051
			y: 0.0
			z: -2.713526
		}, Vertex{
			x: -1.677051
			y: 0.0
			z: 2.713526
		}, Vertex{
			x: -1.677051
			y: 0.0
			z: -2.713526
		}, Vertex{
			x: 2.713526
			y: 1.677051
			z: 0.0
		}, Vertex{
			x: 2.713526
			y: -1.677051
			z: 0.0
		}, Vertex{
			x: -2.713526
			y: 1.677051
			z: 0.0
		}, Vertex{
			x: -2.713526
			y: -1.677051
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 2.713526
			z: 1.677051
		}, Vertex{
			x: 0.0
			y: 2.713526
			z: -1.677051
		}, Vertex{
			x: 0.0
			y: -2.713526
			z: 1.677051
		}, Vertex{
			x: 0.0
			y: -2.713526
			z: -1.677051
		}, Vertex{
			x: 0.0
			y: 0.7725425
			z: 2.022543
		}, Vertex{
			x: 0.0
			y: 0.7725425
			z: -2.022543
		}, Vertex{
			x: 0.0
			y: -0.7725425
			z: 2.022543
		}, Vertex{
			x: 0.0
			y: -0.7725425
			z: -2.022543
		}, Vertex{
			x: 2.022543
			y: 0.0
			z: 0.7725425
		}, Vertex{
			x: 2.022543
			y: 0.0
			z: -0.7725425
		}, Vertex{
			x: -2.022543
			y: 0.0
			z: 0.7725425
		}, Vertex{
			x: -2.022543
			y: 0.0
			z: -0.7725425
		}, Vertex{
			x: 0.7725425
			y: 2.022543
			z: 0.0
		}, Vertex{
			x: 0.7725425
			y: -2.022543
			z: 0.0
		}, Vertex{
			x: -0.7725425
			y: 2.022543
			z: 0.0
		}, Vertex{
			x: -0.7725425
			y: -2.022543
			z: 0.0
		}, Vertex{
			x: 1.036475
			y: 0.0
			z: 1.677051
		}, Vertex{
			x: 1.036475
			y: 0.0
			z: -1.677051
		}, Vertex{
			x: -1.036475
			y: 0.0
			z: 1.677051
		}, Vertex{
			x: -1.036475
			y: 0.0
			z: -1.677051
		}, Vertex{
			x: 1.677051
			y: 1.036475
			z: 0.0
		}, Vertex{
			x: 1.677051
			y: -1.036475
			z: 0.0
		}, Vertex{
			x: -1.677051
			y: 1.036475
			z: 0.0
		}, Vertex{
			x: -1.677051
			y: -1.036475
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.677051
			z: 1.036475
		}, Vertex{
			x: 0.0
			y: 1.677051
			z: -1.036475
		}, Vertex{
			x: 0.0
			y: -1.677051
			z: 1.036475
		}, Vertex{
			x: 0.0
			y: -1.677051
			z: -1.036475
		}, Vertex{
			x: 1.25
			y: 1.25
			z: 1.25
		}, Vertex{
			x: 1.25
			y: 1.25
			z: -1.25
		}, Vertex{
			x: 1.25
			y: -1.25
			z: 1.25
		}, Vertex{
			x: 1.25
			y: -1.25
			z: -1.25
		}, Vertex{
			x: -1.25
			y: 1.25
			z: 1.25
		}, Vertex{
			x: -1.25
			y: 1.25
			z: -1.25
		}, Vertex{
			x: -1.25
			y: -1.25
			z: 1.25
		}, Vertex{
			x: -1.25
			y: -1.25
			z: -1.25
		}]
		faces:     [[0, 17, 28], [0, 28, 20], [0, 20, 32], [0, 32, 40],
			[0, 40, 26], [0, 26, 42], [0, 42, 34], [0, 34, 21],
			[0, 21, 29], [0, 29, 17], [1, 16, 29], [1, 29, 21],
			[1, 21, 35], [1, 35, 43], [1, 43, 27], [1, 27, 41],
			[1, 41, 33], [1, 33, 20], [1, 20, 28], [1, 28, 16],
			[2, 19, 31], [2, 31, 23], [2, 23, 34], [2, 34, 38],
			[2, 38, 24], [2, 24, 36], [2, 36, 32], [2, 32, 22],
			[2, 22, 30], [2, 30, 19], [3, 18, 30], [3, 30, 22],
			[3, 22, 33], [3, 33, 37], [3, 37, 25], [3, 25, 39],
			[3, 39, 35], [3, 35, 23], [3, 23, 31], [3, 31, 18],
			[4, 12, 24], [4, 24, 38], [4, 38, 29], [4, 29, 39],
			[4, 39, 25], [4, 25, 13], [4, 13, 33], [4, 33, 22],
			[4, 22, 32], [4, 32, 12], [5, 14, 34], [5, 34, 23],
			[5, 23, 35], [5, 35, 15], [5, 15, 25], [5, 25, 37],
			[5, 37, 28], [5, 28, 36], [5, 36, 24], [5, 24, 14],
			[6, 12, 32], [6, 32, 20], [6, 20, 33], [6, 33, 13],
			[6, 13, 27], [6, 27, 43], [6, 43, 31], [6, 31, 42],
			[6, 42, 26], [6, 26, 12], [7, 14, 26], [7, 26, 40],
			[7, 40, 30], [7, 30, 41], [7, 41, 27], [7, 27, 15],
			[7, 15, 35], [7, 35, 21], [7, 21, 34], [7, 34, 14],
			[8, 14, 24], [8, 24, 16], [8, 16, 28], [8, 28, 37],
			[8, 37, 33], [8, 33, 41], [8, 41, 30], [8, 30, 18],
			[8, 18, 26], [8, 26, 14], [9, 15, 27], [9, 27, 19],
			[9, 19, 30], [9, 30, 40], [9, 40, 32], [9, 32, 36],
			[9, 36, 28], [9, 28, 17], [9, 17, 25], [9, 25, 15],
			[10, 12, 26], [10, 26, 18], [10, 18, 31], [10, 31, 43],
			[10, 43, 35], [10, 35, 39], [10, 39, 29], [10, 29, 16],
			[10, 16, 24], [10, 24, 12], [11, 13, 25], [11, 25, 17],
			[11, 17, 29], [11, 29, 38], [11, 38, 34], [11, 34, 42],
			[11, 42, 31], [11, 31, 19], [11, 19, 27], [11, 27, 13]]
	},
	Polyhedron{
		name:      'GreatDodecahemidodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 0.618034
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -0.618034
		}, Vertex{
			x: 0.0
			y: 0.618034
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -0.618034
			z: 0.0
		}, Vertex{
			x: 0.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -0.618034
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: -0.1909830
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: 0.1909830
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: -0.1909830
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: 0.1909830
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: -0.1909830
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.1909830
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: 0.1909830
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: 0.1909830
			z: -0.309017
		}, Vertex{
			x: -0.1909830
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: -0.1909830
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: -0.1909830
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: 0.1909830
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: 0.1909830
			y: -0.309017
			z: 0.5
		}]
		faces:     [[0, 6, 22, 23, 7, 1, 13, 29, 28, 12], [0, 8, 24, 25, 9, 1, 11, 27, 26, 10],
			[2, 14, 6, 10, 18, 3, 21, 13, 9, 17], [2, 15, 7, 11, 19, 3, 20, 12, 8, 16],
			[4, 22, 14, 16, 24, 5, 29, 21, 19, 27], [4, 23, 15, 17, 25, 5, 28, 20, 18, 26],
			[0, 8, 16, 14, 6], [0, 10, 18, 20, 12], [1, 7, 15, 17, 9],
			[1, 13, 21, 19, 11], [2, 15, 23, 22, 14], [2, 16, 24, 25, 17],
			[3, 18, 26, 27, 19], [3, 21, 29, 28, 20], [4, 23, 7, 11, 27],
			[4, 26, 10, 6, 22], [5, 24, 8, 12, 28], [5, 29, 13, 9, 25]]
	},
	Polyhedron{
		name:      'GreatDitrigonalDodecacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.927051
			z: -0.572949
		}, Vertex{
			x: 0.0
			y: 0.927051
			z: 0.572949
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: -0.572949
		}, Vertex{
			x: 0.0
			y: -0.927051
			z: 0.572949
		}, Vertex{
			x: 0.927051
			y: -0.572949
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: -0.572949
			z: 0.0
		}, Vertex{
			x: 0.927051
			y: 0.572949
			z: 0.0
		}, Vertex{
			x: -0.927051
			y: 0.572949
			z: 0.0
		}, Vertex{
			x: -0.572949
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: -0.572949
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: 0.572949
			y: 0.0
			z: 0.927051
		}, Vertex{
			x: 0.572949
			y: 0.0
			z: -0.927051
		}, Vertex{
			x: 0.9917610
			y: 0.0
			z: 0.378819
		}, Vertex{
			x: 0.9917610
			y: 0.0
			z: -0.378819
		}, Vertex{
			x: -0.9917610
			y: 0.0
			z: 0.378819
		}, Vertex{
			x: -0.9917610
			y: 0.0
			z: -0.378819
		}, Vertex{
			x: 0.0
			y: 0.378819
			z: 0.9917610
		}, Vertex{
			x: 0.0
			y: 0.378819
			z: -0.9917610
		}, Vertex{
			x: 0.0
			y: -0.378819
			z: 0.9917610
		}, Vertex{
			x: 0.0
			y: -0.378819
			z: -0.9917610
		}, Vertex{
			x: 0.378819
			y: 0.9917610
			z: 0.0
		}, Vertex{
			x: -0.378819
			y: 0.9917610
			z: 0.0
		}, Vertex{
			x: 0.378819
			y: -0.9917610
			z: 0.0
		}, Vertex{
			x: -0.378819
			y: -0.9917610
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.175186
			z: 0.7263052
		}, Vertex{
			x: 0.0
			y: -1.175186
			z: -0.7263052
		}, Vertex{
			x: 0.0
			y: 1.175186
			z: 0.7263052
		}, Vertex{
			x: 0.0
			y: 1.175186
			z: -0.7263052
		}, Vertex{
			x: -1.175186
			y: 0.7263052
			z: 0.0
		}, Vertex{
			x: 1.175186
			y: 0.7263052
			z: 0.0
		}, Vertex{
			x: -1.175186
			y: -0.7263052
			z: 0.0
		}, Vertex{
			x: 1.175186
			y: -0.7263052
			z: 0.0
		}, Vertex{
			x: 0.7263052
			y: 0.0
			z: -1.175186
		}, Vertex{
			x: 0.7263052
			y: 0.0
			z: 1.175186
		}, Vertex{
			x: -0.7263052
			y: 0.0
			z: -1.175186
		}, Vertex{
			x: -0.7263052
			y: 0.0
			z: 1.175186
		}, Vertex{
			x: -0.612942
			y: -0.612942
			z: -0.612942
		}, Vertex{
			x: -0.612942
			y: -0.612942
			z: 0.612942
		}, Vertex{
			x: 0.612942
			y: -0.612942
			z: -0.612942
		}, Vertex{
			x: 0.612942
			y: -0.612942
			z: 0.612942
		}, Vertex{
			x: -0.612942
			y: 0.612942
			z: -0.612942
		}, Vertex{
			x: -0.612942
			y: 0.612942
			z: 0.612942
		}, Vertex{
			x: 0.612942
			y: 0.612942
			z: -0.612942
		}, Vertex{
			x: 0.612942
			y: 0.612942
			z: 0.612942
		}]
		faces:     [[24, 2, 38, 4], [24, 4, 12, 10], [24, 10, 16, 8],
			[24, 8, 14, 5], [24, 5, 36, 2], [25, 4, 39, 3], [25, 3, 37, 5],
			[25, 5, 15, 9], [25, 9, 17, 11], [25, 11, 13, 4],
			[26, 0, 40, 7], [26, 7, 14, 8], [26, 8, 18, 10], [26, 10, 12, 6],
			[26, 6, 42, 0], [27, 1, 43, 6], [27, 6, 13, 11], [27, 11, 19, 9],
			[27, 9, 15, 7], [27, 7, 41, 1], [28, 0, 17, 9], [28, 9, 36, 5],
			[28, 5, 37, 8], [28, 8, 16, 1], [28, 1, 20, 0], [29, 0, 21, 1],
			[29, 1, 16, 10], [29, 10, 39, 4], [29, 4, 38, 11],
			[29, 11, 17, 0], [30, 2, 22, 3], [30, 3, 18, 8], [30, 8, 41, 7],
			[30, 7, 40, 9], [30, 9, 19, 2], [31, 2, 19, 11], [31, 11, 42, 6],
			[31, 6, 43, 10], [31, 10, 18, 3], [31, 3, 23, 2],
			[32, 0, 20, 6], [32, 6, 12, 4], [32, 4, 22, 2], [32, 2, 36, 9],
			[32, 9, 40, 0], [33, 1, 41, 8], [33, 8, 37, 3], [33, 3, 22, 4],
			[33, 4, 13, 6], [33, 6, 20, 1], [34, 0, 42, 11], [34, 11, 38, 2],
			[34, 2, 23, 5], [34, 5, 14, 7], [34, 7, 21, 0], [35, 1, 21, 7],
			[35, 7, 15, 5], [35, 5, 23, 3], [35, 3, 39, 10], [35, 10, 43, 1]]
	},
	Polyhedron{
		name:      'MedialDeltoidalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.341641
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.341641
		}, Vertex{
			x: 1.341641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.341641
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.341641
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.341641
			z: 0.0
		}, Vertex{
			x: 0.7783914
			y: 0.0
			z: 1.259464
		}, Vertex{
			x: 0.7783914
			y: 0.0
			z: -1.259464
		}, Vertex{
			x: -0.7783914
			y: 0.0
			z: 1.259464
		}, Vertex{
			x: -0.7783914
			y: 0.0
			z: -1.259464
		}, Vertex{
			x: 1.259464
			y: 0.7783914
			z: 0.0
		}, Vertex{
			x: 1.259464
			y: -0.7783914
			z: 0.0
		}, Vertex{
			x: -1.259464
			y: 0.7783914
			z: 0.0
		}, Vertex{
			x: -1.259464
			y: -0.7783914
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.259464
			z: 0.7783914
		}, Vertex{
			x: 0.0
			y: 1.259464
			z: -0.7783914
		}, Vertex{
			x: 0.0
			y: -1.259464
			z: 0.7783914
		}, Vertex{
			x: 0.0
			y: -1.259464
			z: -0.7783914
		}, Vertex{
			x: 0.4145898
			y: 0.6708204
			z: 1.085410
		}, Vertex{
			x: 0.4145898
			y: 0.6708204
			z: -1.085410
		}, Vertex{
			x: 0.4145898
			y: -0.6708204
			z: 1.085410
		}, Vertex{
			x: 0.4145898
			y: -0.6708204
			z: -1.085410
		}, Vertex{
			x: -0.4145898
			y: 0.6708204
			z: 1.085410
		}, Vertex{
			x: -0.4145898
			y: 0.6708204
			z: -1.085410
		}, Vertex{
			x: -0.4145898
			y: -0.6708204
			z: 1.085410
		}, Vertex{
			x: -0.4145898
			y: -0.6708204
			z: -1.085410
		}, Vertex{
			x: 1.085410
			y: 0.4145898
			z: 0.6708204
		}, Vertex{
			x: 1.085410
			y: 0.4145898
			z: -0.6708204
		}, Vertex{
			x: 1.085410
			y: -0.4145898
			z: 0.6708204
		}, Vertex{
			x: 1.085410
			y: -0.4145898
			z: -0.6708204
		}, Vertex{
			x: -1.085410
			y: 0.4145898
			z: 0.6708204
		}, Vertex{
			x: -1.085410
			y: 0.4145898
			z: -0.6708204
		}, Vertex{
			x: -1.085410
			y: -0.4145898
			z: 0.6708204
		}, Vertex{
			x: -1.085410
			y: -0.4145898
			z: -0.6708204
		}, Vertex{
			x: 0.6708204
			y: 1.085410
			z: 0.4145898
		}, Vertex{
			x: 0.6708204
			y: 1.085410
			z: -0.4145898
		}, Vertex{
			x: 0.6708204
			y: -1.085410
			z: 0.4145898
		}, Vertex{
			x: 0.6708204
			y: -1.085410
			z: -0.4145898
		}, Vertex{
			x: -0.6708204
			y: 1.085410
			z: 0.4145898
		}, Vertex{
			x: -0.6708204
			y: 1.085410
			z: -0.4145898
		}, Vertex{
			x: -0.6708204
			y: -1.085410
			z: 0.4145898
		}, Vertex{
			x: -0.6708204
			y: -1.085410
			z: -0.4145898
		}, Vertex{
			x: 0.6496271
			y: 0.0
			z: 1.051119
		}, Vertex{
			x: 0.6496271
			y: 0.0
			z: -1.051119
		}, Vertex{
			x: -0.6496271
			y: 0.0
			z: 1.051119
		}, Vertex{
			x: -0.6496271
			y: 0.0
			z: -1.051119
		}, Vertex{
			x: 1.051119
			y: 0.6496271
			z: 0.0
		}, Vertex{
			x: 1.051119
			y: -0.6496271
			z: 0.0
		}, Vertex{
			x: -1.051119
			y: 0.6496271
			z: 0.0
		}, Vertex{
			x: -1.051119
			y: -0.6496271
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.051119
			z: 0.6496271
		}, Vertex{
			x: 0.0
			y: 1.051119
			z: -0.6496271
		}, Vertex{
			x: 0.0
			y: -1.051119
			z: 0.6496271
		}, Vertex{
			x: 0.0
			y: -1.051119
			z: -0.6496271
		}]
		faces:     [[6, 2, 46, 34], [6, 34, 50, 22], [6, 22, 44, 24],
			[6, 24, 52, 36], [6, 36, 47, 2], [7, 2, 47, 37], [7, 37, 53, 25],
			[7, 25, 45, 23], [7, 23, 51, 35], [7, 35, 46, 2],
			[8, 3, 49, 40], [8, 40, 52, 20], [8, 20, 42, 18],
			[8, 18, 50, 38], [8, 38, 48, 3], [9, 3, 48, 39], [9, 39, 51, 19],
			[9, 19, 43, 21], [9, 21, 53, 41], [9, 41, 49, 3],
			[10, 4, 50, 18], [10, 18, 42, 28], [10, 28, 47, 29],
			[10, 29, 43, 19], [10, 19, 51, 4], [11, 5, 53, 21],
			[11, 21, 43, 27], [11, 27, 46, 26], [11, 26, 42, 20],
			[11, 20, 52, 5], [12, 4, 51, 23], [12, 23, 45, 33],
			[12, 33, 49, 32], [12, 32, 44, 22], [12, 22, 50, 4],
			[13, 5, 52, 24], [13, 24, 44, 30], [13, 30, 48, 31],
			[13, 31, 45, 25], [13, 25, 53, 5], [14, 0, 42, 26],
			[14, 26, 46, 35], [14, 35, 51, 39], [14, 39, 48, 30],
			[14, 30, 44, 0], [15, 1, 45, 31], [15, 31, 48, 38],
			[15, 38, 50, 34], [15, 34, 46, 27], [15, 27, 43, 1],
			[16, 0, 44, 32], [16, 32, 49, 41], [16, 41, 53, 37],
			[16, 37, 47, 28], [16, 28, 42, 0], [17, 1, 43, 29],
			[17, 29, 47, 36], [17, 36, 52, 40], [17, 40, 49, 33],
			[17, 33, 45, 1]]
	},
	Polyhedron{
		name:      'MedialHexagonalHexecontahedron'
		vertexes_: [Vertex{
			x: 0.7254514
			y: 0.0
			z: 1.173805
		}, Vertex{
			x: 0.7254514
			y: 0.0
			z: -1.173805
		}, Vertex{
			x: -0.7254514
			y: 0.0
			z: 1.173805
		}, Vertex{
			x: -0.7254514
			y: 0.0
			z: -1.173805
		}, Vertex{
			x: 1.173805
			y: 0.7254514
			z: 0.0
		}, Vertex{
			x: 1.173805
			y: -0.7254514
			z: 0.0
		}, Vertex{
			x: -1.173805
			y: 0.7254514
			z: 0.0
		}, Vertex{
			x: -1.173805
			y: -0.7254514
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.173805
			z: 0.7254514
		}, Vertex{
			x: 0.0
			y: 1.173805
			z: -0.7254514
		}, Vertex{
			x: 0.0
			y: -1.173805
			z: 0.7254514
		}, Vertex{
			x: 0.0
			y: -1.173805
			z: -0.7254514
		}, Vertex{
			x: 0.0
			y: 0.3760450
			z: 0.9844984
		}, Vertex{
			x: 0.0
			y: 0.3760450
			z: -0.9844984
		}, Vertex{
			x: 0.0
			y: -0.3760450
			z: 0.9844984
		}, Vertex{
			x: 0.0
			y: -0.3760450
			z: -0.9844984
		}, Vertex{
			x: 0.9844984
			y: 0.0
			z: 0.3760450
		}, Vertex{
			x: 0.9844984
			y: 0.0
			z: -0.3760450
		}, Vertex{
			x: -0.9844984
			y: 0.0
			z: 0.3760450
		}, Vertex{
			x: -0.9844984
			y: 0.0
			z: -0.3760450
		}, Vertex{
			x: 0.3760450
			y: 0.9844984
			z: 0.0
		}, Vertex{
			x: 0.3760450
			y: -0.9844984
			z: 0.0
		}, Vertex{
			x: -0.3760450
			y: 0.9844984
			z: 0.0
		}, Vertex{
			x: -0.3760450
			y: -0.9844984
			z: 0.0
		}, Vertex{
			x: 0.4388984
			y: 0.03581639
			z: 0.9574615
		}, Vertex{
			x: 0.4388984
			y: -0.03581639
			z: -0.9574615
		}, Vertex{
			x: -0.4388984
			y: -0.03581639
			z: 0.9574615
		}, Vertex{
			x: -0.4388984
			y: 0.03581639
			z: -0.9574615
		}, Vertex{
			x: 0.9574615
			y: 0.4388984
			z: 0.03581639
		}, Vertex{
			x: 0.9574615
			y: -0.4388984
			z: -0.03581639
		}, Vertex{
			x: -0.9574615
			y: -0.4388984
			z: 0.03581639
		}, Vertex{
			x: -0.9574615
			y: 0.4388984
			z: -0.03581639
		}, Vertex{
			x: 0.03581639
			y: 0.9574615
			z: 0.4388984
		}, Vertex{
			x: 0.03581639
			y: -0.9574615
			z: -0.4388984
		}, Vertex{
			x: -0.03581639
			y: -0.9574615
			z: 0.4388984
		}, Vertex{
			x: -0.03581639
			y: 0.9574615
			z: -0.4388984
		}, Vertex{
			x: 0.4863450
			y: -0.1125866
			z: 0.9281378
		}, Vertex{
			x: 0.4863450
			y: 0.1125866
			z: -0.9281378
		}, Vertex{
			x: -0.4863450
			y: 0.1125866
			z: 0.9281378
		}, Vertex{
			x: -0.4863450
			y: -0.1125866
			z: -0.9281378
		}, Vertex{
			x: 0.9281378
			y: -0.4863450
			z: 0.1125866
		}, Vertex{
			x: 0.9281378
			y: 0.4863450
			z: -0.1125866
		}, Vertex{
			x: -0.9281378
			y: 0.4863450
			z: 0.1125866
		}, Vertex{
			x: -0.9281378
			y: -0.4863450
			z: -0.1125866
		}, Vertex{
			x: 0.1125866
			y: -0.9281378
			z: 0.4863450
		}, Vertex{
			x: 0.1125866
			y: 0.9281378
			z: -0.4863450
		}, Vertex{
			x: -0.1125866
			y: 0.9281378
			z: 0.4863450
		}, Vertex{
			x: -0.1125866
			y: -0.9281378
			z: -0.4863450
		}, Vertex{
			x: 0.5442971
			y: 0.1347224
			z: 0.8923215
		}, Vertex{
			x: 0.5442971
			y: -0.1347224
			z: -0.8923215
		}, Vertex{
			x: -0.5442971
			y: -0.1347224
			z: 0.8923215
		}, Vertex{
			x: -0.5442971
			y: 0.1347224
			z: -0.8923215
		}, Vertex{
			x: 0.8923215
			y: 0.5442971
			z: 0.1347224
		}, Vertex{
			x: 0.8923215
			y: -0.5442971
			z: -0.1347224
		}, Vertex{
			x: -0.8923215
			y: -0.5442971
			z: 0.1347224
		}, Vertex{
			x: -0.8923215
			y: 0.5442971
			z: -0.1347224
		}, Vertex{
			x: 0.1347224
			y: 0.8923215
			z: 0.5442971
		}, Vertex{
			x: 0.1347224
			y: -0.8923215
			z: -0.5442971
		}, Vertex{
			x: -0.1347224
			y: -0.8923215
			z: 0.5442971
		}, Vertex{
			x: -0.1347224
			y: 0.8923215
			z: -0.5442971
		}, Vertex{
			x: 0.5379422
			y: 0.0
			z: 0.8704088
		}, Vertex{
			x: 0.5379422
			y: 0.0
			z: -0.8704088
		}, Vertex{
			x: -0.5379422
			y: 0.0
			z: 0.8704088
		}, Vertex{
			x: -0.5379422
			y: 0.0
			z: -0.8704088
		}, Vertex{
			x: 0.8704088
			y: 0.5379422
			z: 0.0
		}, Vertex{
			x: 0.8704088
			y: -0.5379422
			z: 0.0
		}, Vertex{
			x: -0.8704088
			y: 0.5379422
			z: 0.0
		}, Vertex{
			x: -0.8704088
			y: -0.5379422
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.8704088
			z: 0.5379422
		}, Vertex{
			x: 0.0
			y: 0.8704088
			z: -0.5379422
		}, Vertex{
			x: 0.0
			y: -0.8704088
			z: 0.5379422
		}, Vertex{
			x: 0.0
			y: -0.8704088
			z: -0.5379422
		}, Vertex{
			x: 0.6210674
			y: -0.1053988
			z: 0.8448748
		}, Vertex{
			x: 0.6210674
			y: 0.1053988
			z: -0.8448748
		}, Vertex{
			x: -0.6210674
			y: 0.1053988
			z: 0.8448748
		}, Vertex{
			x: -0.6210674
			y: -0.1053988
			z: -0.8448748
		}, Vertex{
			x: 0.8448748
			y: -0.6210674
			z: 0.1053988
		}, Vertex{
			x: 0.8448748
			y: 0.6210674
			z: -0.1053988
		}, Vertex{
			x: -0.8448748
			y: 0.6210674
			z: 0.1053988
		}, Vertex{
			x: -0.8448748
			y: -0.6210674
			z: -0.1053988
		}, Vertex{
			x: 0.1053988
			y: -0.8448748
			z: 0.6210674
		}, Vertex{
			x: 0.1053988
			y: 0.8448748
			z: -0.6210674
		}, Vertex{
			x: -0.1053988
			y: 0.8448748
			z: 0.6210674
		}, Vertex{
			x: -0.1053988
			y: -0.8448748
			z: -0.6210674
		}, Vertex{
			x: 0.6568838
			y: 0.04744662
			z: 0.8227391
		}, Vertex{
			x: 0.6568838
			y: -0.04744662
			z: -0.8227391
		}, Vertex{
			x: -0.6568838
			y: -0.04744662
			z: 0.8227391
		}, Vertex{
			x: -0.6568838
			y: 0.04744662
			z: -0.8227391
		}, Vertex{
			x: 0.8227391
			y: 0.6568838
			z: 0.04744662
		}, Vertex{
			x: 0.8227391
			y: -0.6568838
			z: -0.04744662
		}, Vertex{
			x: -0.8227391
			y: -0.6568838
			z: 0.04744662
		}, Vertex{
			x: -0.8227391
			y: 0.6568838
			z: -0.04744662
		}, Vertex{
			x: 0.04744662
			y: 0.8227391
			z: 0.6568838
		}, Vertex{
			x: 0.04744662
			y: -0.8227391
			z: -0.6568838
		}, Vertex{
			x: -0.04744662
			y: -0.8227391
			z: 0.6568838
		}, Vertex{
			x: -0.04744662
			y: 0.8227391
			z: -0.6568838
		}, Vertex{
			x: 0.6084535
			y: 0.6084535
			z: 0.6084535
		}, Vertex{
			x: 0.6084535
			y: 0.6084535
			z: -0.6084535
		}, Vertex{
			x: 0.6084535
			y: -0.6084535
			z: 0.6084535
		}, Vertex{
			x: 0.6084535
			y: -0.6084535
			z: -0.6084535
		}, Vertex{
			x: -0.6084535
			y: 0.6084535
			z: 0.6084535
		}, Vertex{
			x: -0.6084535
			y: 0.6084535
			z: -0.6084535
		}, Vertex{
			x: -0.6084535
			y: -0.6084535
			z: 0.6084535
		}, Vertex{
			x: -0.6084535
			y: -0.6084535
			z: -0.6084535
		}]
		faces:     [[0, 28, 64, 77, 20, 56], [0, 56, 68, 46, 100, 38],
			[0, 38, 62, 86, 102, 94], [0, 94, 70, 34, 21, 76],
			[0, 76, 65, 53, 17, 28], [1, 29, 65, 76, 21, 57],
			[1, 57, 71, 47, 103, 39], [1, 39, 63, 87, 101, 95],
			[1, 95, 69, 35, 20, 77], [1, 77, 64, 52, 16, 29],
			[2, 30, 67, 79, 23, 58], [2, 58, 70, 44, 98, 36],
			[2, 36, 60, 84, 96, 92], [2, 92, 68, 32, 22, 78],
			[2, 78, 66, 55, 19, 30], [3, 31, 66, 78, 22, 59],
			[3, 59, 69, 45, 97, 37], [3, 37, 61, 85, 99, 93],
			[3, 93, 71, 33, 23, 79], [3, 79, 67, 54, 18, 31],
			[4, 32, 68, 82, 12, 48], [4, 48, 60, 36, 98, 40],
			[4, 40, 65, 89, 99, 85], [4, 85, 61, 25, 13, 81],
			[4, 81, 69, 59, 22, 32], [5, 33, 71, 83, 15, 49],
			[5, 49, 61, 37, 97, 41], [5, 41, 64, 88, 96, 84],
			[5, 84, 60, 24, 14, 80], [5, 80, 70, 58, 23, 33],
			[6, 35, 69, 81, 13, 51], [6, 51, 63, 39, 103, 43],
			[6, 43, 67, 90, 102, 86], [6, 86, 62, 26, 12, 82],
			[6, 82, 68, 56, 20, 35], [7, 34, 70, 80, 14, 50],
			[7, 50, 62, 38, 100, 42], [7, 42, 66, 91, 101, 87],
			[7, 87, 63, 27, 15, 83], [7, 83, 71, 57, 21, 34],
			[8, 24, 60, 72, 16, 52], [8, 52, 64, 41, 97, 45],
			[8, 45, 69, 95, 101, 91], [8, 91, 66, 31, 18, 74],
			[8, 74, 62, 50, 14, 24], [9, 27, 63, 75, 19, 55],
			[9, 55, 66, 42, 100, 46], [9, 46, 68, 92, 96, 88],
			[9, 88, 64, 28, 17, 73], [9, 73, 61, 49, 15, 27],
			[10, 26, 62, 74, 18, 54], [10, 54, 67, 43, 103, 47],
			[10, 47, 71, 93, 99, 89], [10, 89, 65, 29, 16, 72],
			[10, 72, 60, 48, 12, 26], [11, 25, 61, 73, 17, 53],
			[11, 53, 65, 40, 98, 44], [11, 44, 70, 94, 102, 90],
			[11, 90, 67, 30, 19, 75], [11, 75, 63, 51, 13, 25]]
	},
	Polyhedron{
		name:      'Rhombicosahedron'
		vertexes_: [Vertex{
			x: 0.1909830
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: 0.1909830
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: 1.309017
		}, Vertex{
			x: -0.1909830
			y: 0.0
			z: -1.309017
		}, Vertex{
			x: 1.309017
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: 1.309017
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: 0.1909830
			z: 0.0
		}, Vertex{
			x: -1.309017
			y: -0.1909830
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: 1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: 0.1909830
		}, Vertex{
			x: 0.0
			y: -1.309017
			z: -0.1909830
		}, Vertex{
			x: 0.5
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: 0.5
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: 0.5
			z: -1.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: 1.118034
		}, Vertex{
			x: -0.5
			y: -0.5
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: 1.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: 0.5
			z: -0.5
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: 0.5
		}, Vertex{
			x: -1.118034
			y: -0.5
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: 0.5
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: 1.118034
			z: -0.5
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: 0.5
		}, Vertex{
			x: -0.5
			y: -1.118034
			z: -0.5
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: 1.0
		}, Vertex{
			x: 0.309017
			y: 0.809017
			z: -1.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: 1.0
		}, Vertex{
			x: 0.309017
			y: -0.809017
			z: -1.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: 1.0
		}, Vertex{
			x: -0.309017
			y: 0.809017
			z: -1.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: 1.0
		}, Vertex{
			x: -0.309017
			y: -0.809017
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: 1.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: 1.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: 1.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: -1.0
			y: 0.309017
			z: 0.809017
		}, Vertex{
			x: -1.0
			y: 0.309017
			z: -0.809017
		}, Vertex{
			x: -1.0
			y: -0.309017
			z: 0.809017
		}, Vertex{
			x: -1.0
			y: -0.309017
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 1.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: 1.0
			z: -0.309017
		}, Vertex{
			x: 0.809017
			y: -1.0
			z: 0.309017
		}, Vertex{
			x: 0.809017
			y: -1.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: 1.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: 1.0
			z: -0.309017
		}, Vertex{
			x: -0.809017
			y: -1.0
			z: 0.309017
		}, Vertex{
			x: -0.809017
			y: -1.0
			z: -0.309017
		}]
		faces:     [[0, 42, 10, 55, 5, 44], [0, 46, 4, 53, 8, 40],
			[2, 36, 8, 57, 6, 50], [2, 48, 7, 59, 10, 38], [15, 13, 53, 20, 22, 55],
			[15, 19, 49, 33, 29, 45], [17, 13, 47, 31, 35, 51],
			[17, 19, 59, 26, 24, 57], [30, 46, 12, 16, 50, 34],
			[30, 42, 26, 27, 43, 31], [32, 48, 18, 14, 44, 28],
			[32, 36, 20, 21, 37, 33], [39, 23, 22, 38, 34, 35],
			[39, 11, 58, 7, 49, 3], [41, 25, 24, 40, 28, 29],
			[41, 9, 52, 4, 47, 1], [54, 11, 43, 1, 45, 5], [54, 23, 21, 52, 12, 14],
			[56, 9, 37, 3, 51, 6], [56, 25, 27, 58, 18, 16], [0, 42, 30, 46],
			[0, 44, 28, 40], [1, 41, 29, 45], [1, 47, 31, 43],
			[3, 39, 35, 51], [3, 49, 33, 37], [5, 44, 14, 54],
			[5, 55, 15, 45], [6, 50, 16, 56], [6, 57, 17, 51],
			[7, 49, 19, 59], [7, 58, 18, 48], [8, 36, 20, 53],
			[8, 57, 24, 40], [9, 41, 25, 56], [9, 52, 21, 37],
			[11, 39, 23, 54], [11, 58, 27, 43], [12, 16, 18, 14],
			[12, 46, 4, 52], [13, 15, 19, 17], [13, 53, 4, 47],
			[22, 23, 21, 20], [22, 38, 10, 55], [26, 24, 25, 27],
			[26, 59, 10, 42], [32, 28, 29, 33], [32, 48, 2, 36],
			[34, 35, 31, 30], [34, 38, 2, 50]]
	},
	Polyhedron{
		name:      'Dodecadodecahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 1.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.0
		}, Vertex{
			x: 1.0
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.0
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.0
			z: 0.0
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: 0.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: 0.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: 0.5
			z: -0.809017
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: 0.809017
		}, Vertex{
			x: -0.309017
			y: -0.5
			z: -0.809017
		}, Vertex{
			x: 0.809017
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: 0.809017
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: 0.809017
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: 0.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: 0.309017
			z: -0.5
		}, Vertex{
			x: -0.809017
			y: -0.309017
			z: 0.5
		}, Vertex{
			x: -0.809017
			y: -0.309017
			z: -0.5
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: 0.809017
			z: -0.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: 0.309017
		}, Vertex{
			x: 0.5
			y: -0.809017
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: 0.809017
			z: -0.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: 0.309017
		}, Vertex{
			x: -0.5
			y: -0.809017
			z: -0.309017
		}]
		faces:     [[0, 14, 23, 27, 18], [0, 18, 12, 10, 20],
			[0, 20, 29, 25, 16], [0, 16, 6, 8, 14], [1, 17, 24, 28, 21],
			[1, 21, 11, 13, 19], [1, 19, 26, 22, 15], [1, 15, 9, 7, 17],
			[2, 22, 10, 12, 24], [2, 24, 17, 16, 25], [2, 25, 13, 11, 23],
			[2, 23, 14, 15, 22], [3, 27, 7, 9, 29], [3, 29, 20, 21, 28],
			[3, 28, 8, 6, 26], [3, 26, 19, 18, 27], [4, 6, 16, 17, 7],
			[4, 7, 27, 23, 11], [4, 11, 21, 20, 10], [4, 10, 22, 26, 6],
			[5, 8, 28, 24, 12], [5, 12, 18, 19, 13], [5, 13, 25, 29, 9],
			[5, 9, 15, 14, 8]]
	},
	Polyhedron{
		name:      'GreatIcosacronicHexecontahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: 0.690983
			z: -1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: 1.809017
		}, Vertex{
			x: 0.0
			y: -0.690983
			z: -1.809017
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: 1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: 0.690983
		}, Vertex{
			x: -1.809017
			y: 0.0
			z: -0.690983
		}, Vertex{
			x: 0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: 0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: 1.809017
			z: 0.0
		}, Vertex{
			x: -0.690983
			y: -1.809017
			z: 0.0
		}, Vertex{
			x: 0.7263052
			y: 0.0
			z: 1.175186
		}, Vertex{
			x: 0.7263052
			y: 0.0
			z: -1.175186
		}, Vertex{
			x: -0.7263052
			y: 0.0
			z: 1.175186
		}, Vertex{
			x: -0.7263052
			y: 0.0
			z: -1.175186
		}, Vertex{
			x: 1.175186
			y: 0.7263052
			z: 0.0
		}, Vertex{
			x: 1.175186
			y: -0.7263052
			z: 0.0
		}, Vertex{
			x: -1.175186
			y: 0.7263052
			z: 0.0
		}, Vertex{
			x: -1.175186
			y: -0.7263052
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.175186
			z: 0.7263052
		}, Vertex{
			x: 0.0
			y: 1.175186
			z: -0.7263052
		}, Vertex{
			x: 0.0
			y: -1.175186
			z: 0.7263052
		}, Vertex{
			x: 0.0
			y: -1.175186
			z: -0.7263052
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: 1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: 1.118034
			z: -1.118034
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: 1.118034
		}, Vertex{
			x: -1.118034
			y: -1.118034
			z: -1.118034
		}, Vertex{
			x: 0.0
			y: 0.378819
			z: 0.9917610
		}, Vertex{
			x: 0.0
			y: 0.378819
			z: -0.9917610
		}, Vertex{
			x: 0.0
			y: -0.378819
			z: 0.9917610
		}, Vertex{
			x: 0.0
			y: -0.378819
			z: -0.9917610
		}, Vertex{
			x: 0.9917610
			y: 0.0
			z: 0.378819
		}, Vertex{
			x: 0.9917610
			y: 0.0
			z: -0.378819
		}, Vertex{
			x: -0.9917610
			y: 0.0
			z: 0.378819
		}, Vertex{
			x: -0.9917610
			y: 0.0
			z: -0.378819
		}, Vertex{
			x: 0.378819
			y: 0.9917610
			z: 0.0
		}, Vertex{
			x: 0.378819
			y: -0.9917610
			z: 0.0
		}, Vertex{
			x: -0.378819
			y: 0.9917610
			z: 0.0
		}, Vertex{
			x: -0.378819
			y: -0.9917610
			z: 0.0
		}, Vertex{
			x: 0.612942
			y: 0.612942
			z: 0.612942
		}, Vertex{
			x: 0.612942
			y: 0.612942
			z: -0.612942
		}, Vertex{
			x: 0.612942
			y: -0.612942
			z: 0.612942
		}, Vertex{
			x: 0.612942
			y: -0.612942
			z: -0.612942
		}, Vertex{
			x: -0.612942
			y: 0.612942
			z: 0.612942
		}, Vertex{
			x: -0.612942
			y: 0.612942
			z: -0.612942
		}, Vertex{
			x: -0.612942
			y: -0.612942
			z: 0.612942
		}, Vertex{
			x: -0.612942
			y: -0.612942
			z: -0.612942
		}]
		faces:     [[12, 6, 50, 11], [12, 11, 41, 27], [12, 27, 37, 25],
			[12, 25, 40, 10], [12, 10, 48, 6], [13, 7, 49, 10],
			[13, 10, 40, 24], [13, 24, 36, 26], [13, 26, 41, 11],
			[13, 11, 51, 7], [14, 4, 44, 8], [14, 8, 42, 29],
			[14, 29, 39, 31], [14, 31, 43, 9], [14, 9, 46, 4],
			[15, 5, 47, 9], [15, 9, 43, 30], [15, 30, 38, 28],
			[15, 28, 42, 8], [15, 8, 45, 5], [16, 2, 46, 9], [16, 9, 47, 3],
			[16, 3, 33, 29], [16, 29, 42, 28], [16, 28, 32, 2],
			[17, 0, 34, 30], [17, 30, 43, 31], [17, 31, 35, 1],
			[17, 1, 45, 8], [17, 8, 44, 0], [18, 2, 32, 24], [18, 24, 40, 25],
			[18, 25, 33, 3], [18, 3, 51, 11], [18, 11, 50, 2],
			[19, 0, 48, 10], [19, 10, 49, 1], [19, 1, 35, 27],
			[19, 27, 41, 26], [19, 26, 34, 0], [20, 1, 49, 7],
			[20, 7, 38, 30], [20, 30, 34, 26], [20, 26, 36, 5],
			[20, 5, 45, 1], [21, 0, 44, 4], [21, 4, 37, 27], [21, 27, 35, 31],
			[21, 31, 39, 6], [21, 6, 48, 0], [22, 3, 47, 5], [22, 5, 36, 24],
			[22, 24, 32, 28], [22, 28, 38, 7], [22, 7, 51, 3],
			[23, 2, 50, 6], [23, 6, 39, 29], [23, 29, 33, 25],
			[23, 25, 37, 4], [23, 4, 46, 2]]
	},
	Polyhedron{
		name:      'PentagonalHexecontahedron(dextro}'
		vertexes_: [Vertex{
			x: 0.1928937
			y: 0.2184834
			z: 2.097054
		}, Vertex{
			x: 0.1928937
			y: -0.2184834
			z: -2.097054
		}, Vertex{
			x: -0.1928937
			y: -0.2184834
			z: 2.097054
		}, Vertex{
			x: -0.1928937
			y: 0.2184834
			z: -2.097054
		}, Vertex{
			x: 2.097054
			y: 0.1928937
			z: 0.2184834
		}, Vertex{
			x: 2.097054
			y: -0.1928937
			z: -0.2184834
		}, Vertex{
			x: -2.097054
			y: -0.1928937
			z: 0.2184834
		}, Vertex{
			x: -2.097054
			y: 0.1928937
			z: -0.2184834
		}, Vertex{
			x: 0.2184834
			y: 2.097054
			z: 0.1928937
		}, Vertex{
			x: 0.2184834
			y: -2.097054
			z: -0.1928937
		}, Vertex{
			x: -0.2184834
			y: -2.097054
			z: 0.1928937
		}, Vertex{
			x: -0.2184834
			y: 2.097054
			z: -0.1928937
		}, Vertex{
			x: 0.0
			y: 0.7554672
			z: 1.977839
		}, Vertex{
			x: 0.0
			y: 0.7554672
			z: -1.977839
		}, Vertex{
			x: 0.0
			y: -0.7554672
			z: 1.977839
		}, Vertex{
			x: 0.0
			y: -0.7554672
			z: -1.977839
		}, Vertex{
			x: 1.977839
			y: 0.0
			z: 0.7554672
		}, Vertex{
			x: 1.977839
			y: 0.0
			z: -0.7554672
		}, Vertex{
			x: -1.977839
			y: 0.0
			z: 0.7554672
		}, Vertex{
			x: -1.977839
			y: 0.0
			z: -0.7554672
		}, Vertex{
			x: 0.7554672
			y: 1.977839
			z: 0.0
		}, Vertex{
			x: 0.7554672
			y: -1.977839
			z: 0.0
		}, Vertex{
			x: -0.7554672
			y: 1.977839
			z: 0.0
		}, Vertex{
			x: -0.7554672
			y: -1.977839
			z: 0.0
		}, Vertex{
			x: 1.167123
			y: 0.0
			z: 1.888445
		}, Vertex{
			x: 1.167123
			y: 0.0
			z: -1.888445
		}, Vertex{
			x: -1.167123
			y: 0.0
			z: 1.888445
		}, Vertex{
			x: -1.167123
			y: 0.0
			z: -1.888445
		}, Vertex{
			x: 1.888445
			y: 1.167123
			z: 0.0
		}, Vertex{
			x: 1.888445
			y: -1.167123
			z: 0.0
		}, Vertex{
			x: -1.888445
			y: 1.167123
			z: 0.0
		}, Vertex{
			x: -1.888445
			y: -1.167123
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.888445
			z: 1.167123
		}, Vertex{
			x: 0.0
			y: 1.888445
			z: -1.167123
		}, Vertex{
			x: 0.0
			y: -1.888445
			z: 1.167123
		}, Vertex{
			x: 0.0
			y: -1.888445
			z: -1.167123
		}, Vertex{
			x: 0.5677154
			y: -0.8249576
			z: 1.865401
		}, Vertex{
			x: 0.5677154
			y: 0.8249576
			z: -1.865401
		}, Vertex{
			x: -0.5677154
			y: 0.8249576
			z: 1.865401
		}, Vertex{
			x: -0.5677154
			y: -0.8249576
			z: -1.865401
		}, Vertex{
			x: 1.865401
			y: -0.5677154
			z: 0.8249576
		}, Vertex{
			x: 1.865401
			y: 0.5677154
			z: -0.8249576
		}, Vertex{
			x: -1.865401
			y: 0.5677154
			z: 0.8249576
		}, Vertex{
			x: -1.865401
			y: -0.5677154
			z: -0.8249576
		}, Vertex{
			x: 0.8249576
			y: -1.865401
			z: 0.5677154
		}, Vertex{
			x: 0.8249576
			y: 1.865401
			z: -0.5677154
		}, Vertex{
			x: -0.8249576
			y: 1.865401
			z: 0.5677154
		}, Vertex{
			x: -0.8249576
			y: -1.865401
			z: -0.5677154
		}, Vertex{
			x: 0.3748217
			y: 1.137066
			z: 1.746187
		}, Vertex{
			x: 0.3748217
			y: -1.137066
			z: -1.746187
		}, Vertex{
			x: -0.3748217
			y: -1.137066
			z: 1.746187
		}, Vertex{
			x: -0.3748217
			y: 1.137066
			z: -1.746187
		}, Vertex{
			x: 1.746187
			y: 0.3748217
			z: 1.137066
		}, Vertex{
			x: 1.746187
			y: -0.3748217
			z: -1.137066
		}, Vertex{
			x: -1.746187
			y: -0.3748217
			z: 1.137066
		}, Vertex{
			x: -1.746187
			y: 0.3748217
			z: -1.137066
		}, Vertex{
			x: 1.137066
			y: 1.746187
			z: 0.3748217
		}, Vertex{
			x: 1.137066
			y: -1.746187
			z: -0.3748217
		}, Vertex{
			x: -1.137066
			y: -1.746187
			z: 0.3748217
		}, Vertex{
			x: -1.137066
			y: 1.746187
			z: -0.3748217
		}, Vertex{
			x: 0.9212289
			y: 0.9599877
			z: 1.646918
		}, Vertex{
			x: 0.9212289
			y: -0.9599877
			z: -1.646918
		}, Vertex{
			x: -0.9212289
			y: -0.9599877
			z: 1.646918
		}, Vertex{
			x: -0.9212289
			y: 0.9599877
			z: -1.646918
		}, Vertex{
			x: 1.646918
			y: 0.9212289
			z: 0.9599877
		}, Vertex{
			x: 1.646918
			y: -0.9212289
			z: -0.9599877
		}, Vertex{
			x: -1.646918
			y: -0.9212289
			z: 0.9599877
		}, Vertex{
			x: -1.646918
			y: 0.9212289
			z: -0.9599877
		}, Vertex{
			x: 0.9599877
			y: 1.646918
			z: 0.9212289
		}, Vertex{
			x: 0.9599877
			y: -1.646918
			z: -0.9212289
		}, Vertex{
			x: -0.9599877
			y: -1.646918
			z: 0.9212289
		}, Vertex{
			x: -0.9599877
			y: 1.646918
			z: -0.9212289
		}, Vertex{
			x: 0.7283352
			y: -1.272096
			z: 1.527703
		}, Vertex{
			x: 0.7283352
			y: 1.272096
			z: -1.527703
		}, Vertex{
			x: -0.7283352
			y: 1.272096
			z: 1.527703
		}, Vertex{
			x: -0.7283352
			y: -1.272096
			z: -1.527703
		}, Vertex{
			x: 1.527703
			y: -0.7283352
			z: 1.272096
		}, Vertex{
			x: 1.527703
			y: 0.7283352
			z: -1.272096
		}, Vertex{
			x: -1.527703
			y: 0.7283352
			z: 1.272096
		}, Vertex{
			x: -1.527703
			y: -0.7283352
			z: -1.272096
		}, Vertex{
			x: 1.272096
			y: -1.527703
			z: 0.7283352
		}, Vertex{
			x: 1.272096
			y: 1.527703
			z: -0.7283352
		}, Vertex{
			x: -1.272096
			y: 1.527703
			z: 0.7283352
		}, Vertex{
			x: -1.272096
			y: -1.527703
			z: -0.7283352
		}, Vertex{
			x: 1.222372
			y: 1.222372
			z: 1.222372
		}, Vertex{
			x: 1.222372
			y: 1.222372
			z: -1.222372
		}, Vertex{
			x: 1.222372
			y: -1.222372
			z: 1.222372
		}, Vertex{
			x: 1.222372
			y: -1.222372
			z: -1.222372
		}, Vertex{
			x: -1.222372
			y: 1.222372
			z: 1.222372
		}, Vertex{
			x: -1.222372
			y: 1.222372
			z: -1.222372
		}, Vertex{
			x: -1.222372
			y: -1.222372
			z: 1.222372
		}, Vertex{
			x: -1.222372
			y: -1.222372
			z: -1.222372
		}]
		faces:     [[24, 0, 2, 14, 36], [24, 36, 72, 86, 76],
			[24, 76, 40, 16, 52], [24, 52, 64, 84, 60], [24, 60, 48, 12, 0],
			[25, 1, 3, 13, 37], [25, 37, 73, 85, 77], [25, 77, 41, 17, 53],
			[25, 53, 65, 87, 61], [25, 61, 49, 15, 1], [26, 2, 0, 12, 38],
			[26, 38, 74, 88, 78], [26, 78, 42, 18, 54], [26, 54, 66, 90, 62],
			[26, 62, 50, 14, 2], [27, 3, 1, 15, 39], [27, 39, 75, 91, 79],
			[27, 79, 43, 19, 55], [27, 55, 67, 89, 63], [27, 63, 51, 13, 3],
			[28, 4, 5, 17, 41], [28, 41, 77, 85, 81], [28, 81, 45, 20, 56],
			[28, 56, 68, 84, 64], [28, 64, 52, 16, 4], [29, 5, 4, 16, 40],
			[29, 40, 76, 86, 80], [29, 80, 44, 21, 57], [29, 57, 69, 87, 65],
			[29, 65, 53, 17, 5], [30, 7, 6, 18, 42], [30, 42, 78, 88, 82],
			[30, 82, 46, 22, 59], [30, 59, 71, 89, 67], [30, 67, 55, 19, 7],
			[31, 6, 7, 19, 43], [31, 43, 79, 91, 83], [31, 83, 47, 23, 58],
			[31, 58, 70, 90, 66], [31, 66, 54, 18, 6], [32, 8, 11, 22, 46],
			[32, 46, 82, 88, 74], [32, 74, 38, 12, 48], [32, 48, 60, 84, 68],
			[32, 68, 56, 20, 8], [33, 11, 8, 20, 45], [33, 45, 81, 85, 73],
			[33, 73, 37, 13, 51], [33, 51, 63, 89, 71], [33, 71, 59, 22, 11],
			[34, 10, 9, 21, 44], [34, 44, 80, 86, 72], [34, 72, 36, 14, 50],
			[34, 50, 62, 90, 70], [34, 70, 58, 23, 10], [35, 9, 10, 23, 47],
			[35, 47, 83, 91, 75], [35, 75, 39, 15, 49], [35, 49, 61, 87, 69],
			[35, 69, 57, 21, 9]]
	},
	Polyhedron{
		name:      'SmallHexacronicIcositetrahedron'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: 3.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -3.414214
		}, Vertex{
			x: 3.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -3.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 3.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -3.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.414214
		}, Vertex{
			x: 0.0
			y: 0.0
			z: -1.414214
		}, Vertex{
			x: 1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: -1.414214
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.414214
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.414214
			z: 0.0
		}, Vertex{
			x: 0.7734591
			y: 0.7734591
			z: 0.7734591
		}, Vertex{
			x: 0.7734591
			y: 0.7734591
			z: -0.7734591
		}, Vertex{
			x: 0.7734591
			y: -0.7734591
			z: 0.7734591
		}, Vertex{
			x: 0.7734591
			y: -0.7734591
			z: -0.7734591
		}, Vertex{
			x: -0.7734591
			y: 0.7734591
			z: 0.7734591
		}, Vertex{
			x: -0.7734591
			y: 0.7734591
			z: -0.7734591
		}, Vertex{
			x: -0.7734591
			y: -0.7734591
			z: 0.7734591
		}, Vertex{
			x: -0.7734591
			y: -0.7734591
			z: -0.7734591
		}]
		faces:     [[12, 0, 8, 4], [12, 4, 6, 2], [12, 2, 10, 0],
			[13, 1, 10, 2], [13, 2, 7, 4], [13, 4, 8, 1], [14, 0, 11, 2],
			[14, 2, 6, 5], [14, 5, 8, 0], [15, 1, 8, 5], [15, 5, 7, 2],
			[15, 2, 11, 1], [16, 0, 10, 3], [16, 3, 6, 4], [16, 4, 9, 0],
			[17, 1, 9, 4], [17, 4, 7, 3], [17, 3, 10, 1], [18, 0, 9, 5],
			[18, 5, 6, 3], [18, 3, 11, 0], [19, 1, 11, 3], [19, 3, 7, 5],
			[19, 5, 9, 1]]
	},
	Polyhedron{
		name:      'PentagonalIcositetrahedron(laevo}'
		vertexes_: [Vertex{
			x: 0.0
			y: 0.0
			z: -1.361410
		}, Vertex{
			x: 0.0
			y: 0.0
			z: 1.361410
		}, Vertex{
			x: -1.361410
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 1.361410
			y: 0.0
			z: 0.0
		}, Vertex{
			x: 0.0
			y: -1.361410
			z: 0.0
		}, Vertex{
			x: 0.0
			y: 1.361410
			z: 0.0
		}, Vertex{
			x: -0.7401838
			y: 0.2187966
			z: -1.023656
		}, Vertex{
			x: -0.7401838
			y: -0.2187966
			z: 1.023656
		}, Vertex{
			x: 0.7401838
			y: -0.2187966
			z: -1.023656
		}, Vertex{
			x: 0.7401838
			y: 0.2187966
			z: 1.023656
		}, Vertex{
			x: -1.023656
			y: 0.7401838
			z: -0.2187966
		}, Vertex{
			x: -1.023656
			y: -0.7401838
			z: 0.2187966
		}, Vertex{
			x: 1.023656
			y: -0.7401838
			z: -0.2187966
		}, Vertex{
			x: 1.023656
			y: 0.7401838
			z: 0.2187966
		}, Vertex{
			x: -0.2187966
			y: 1.023656
			z: -0.7401838
		}, Vertex{
			x: -0.2187966
			y: -1.023656
			z: 0.7401838
		}, Vertex{
			x: 0.2187966
			y: -1.023656
			z: -0.7401838
		}, Vertex{
			x: 0.2187966
			y: 1.023656
			z: 0.7401838
		}, Vertex{
			x: -0.2187966
			y: -0.7401838
			z: -1.023656
		}, Vertex{
			x: -0.2187966
			y: 0.7401838
			z: 1.023656
		}, Vertex{
			x: 0.2187966
			y: 0.7401838
			z: -1.023656
		}, Vertex{
			x: 0.2187966
			y: -0.7401838
			z: 1.023656
		}, Vertex{
			x: -1.023656
			y: -0.2187966
			z: -0.7401838
		}, Vertex{
			x: -1.023656
			y: 0.2187966
			z: 0.7401838
		}, Vertex{
			x: 1.023656
			y: 0.2187966
			z: -0.7401838
		}, Vertex{
			x: 1.023656
			y: -0.2187966
			z: 0.7401838
		}, Vertex{
			x: -0.7401838
			y: -1.023656
			z: -0.2187966
		}, Vertex{
			x: -0.7401838
			y: 1.023656
			z: 0.2187966
		}, Vertex{
			x: 0.7401838
			y: 1.023656
			z: -0.2187966
		}, Vertex{
			x: 0.7401838
			y: -1.023656
			z: 0.2187966
		}, Vertex{
			x: -0.7401838
			y: -0.7401838
			z: -0.7401838
		}, Vertex{
			x: -0.7401838
			y: -0.7401838
			z: 0.7401838
		}, Vertex{
			x: -0.7401838
			y: 0.7401838
			z: -0.7401838
		}, Vertex{
			x: -0.7401838
			y: 0.7401838
			z: 0.7401838
		}, Vertex{
			x: 0.7401838
			y: -0.7401838
			z: -0.7401838
		}, Vertex{
			x: 0.7401838
			y: -0.7401838
			z: 0.7401838
		}, Vertex{
			x: 0.7401838
			y: 0.7401838
			z: -0.7401838
		}, Vertex{
			x: 0.7401838
			y: 0.7401838
			z: 0.7401838
		}]
		faces:     [[0, 18, 30, 22, 6], [0, 8, 34, 16, 18], [0, 20, 36, 24, 8],
			[0, 6, 32, 14, 20], [1, 19, 33, 23, 7], [1, 9, 37, 17, 19],
			[1, 21, 35, 25, 9], [1, 7, 31, 15, 21], [2, 23, 33, 27, 10],
			[2, 11, 31, 7, 23], [2, 22, 30, 26, 11], [2, 10, 32, 6, 22],
			[3, 25, 35, 29, 12], [3, 13, 37, 9, 25], [3, 24, 36, 28, 13],
			[3, 12, 34, 8, 24], [4, 29, 35, 21, 15], [4, 16, 34, 12, 29],
			[4, 26, 30, 18, 16], [4, 15, 31, 11, 26], [5, 28, 36, 20, 14],
			[5, 17, 37, 13, 28], [5, 27, 33, 19, 17], [5, 14, 32, 10, 27]]
	},
]
