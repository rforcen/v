module main

import voronoi


fn ui_obj() {
	voronoi.ui_glfw()
}

fn main() {
	ui_obj()
}
