module main

import queens { gui }

fn main() {
	gui()
}
