module main

import numv as nv { test01, test02, test03, test04, test05, test06, test07, test08 }

fn main() {
	// test01()
	// test02()
	// test03()
	// test04()
	// test05()
	//test06()
	// test07()
	test08()
}
