// johnson polys 1..92

module poly

pub const johnson = [
	&Polyhedron{
		name:     'j1'
		vertexes: [[f32(-0.729665), f32(0.670121), f32(0.319155)],
			[f32(-0.655235), f32(-0.29213), f32(-0.754096)],
			[f32(-0.093922), f32(-0.607123),
				f32(0.537818)],
			[f32(0.702196), f32(0.595691), f32(0.485187)],
			[f32(0.776626), f32(-0.36656),
				f32(-0.588064)]]
		faces:    [[1, 4, 2], [0, 1, 2], [3, 0, 2], [4, 3, 2],
			[4, 1, 0, 3]]
	},
	&Polyhedron{
		name:     'j2'
		vertexes: [[f32(-0.868849), f32(-0.100041), f32(0.61257)],
			[f32(-0.329458), f32(0.976099), f32(0.28078)],
			[f32(-0.26629), f32(-0.013796),
				f32(-0.477654)],
			[f32(-0.13392), f32(-1.03411), f32(0.229829)],
			[f32(0.738834), f32(0.707117),
				f32(-0.307018)],
			[f32(0.859683), f32(-0.535264), f32(-0.338508)]]
		faces:    [[3, 0, 2], [5, 3, 2], [4, 5, 2], [1, 4, 2],
			[0, 1, 2], [0, 3, 5, 4, 1]]
	},
	&Polyhedron{
		name:     'j3'
		vertexes: [[f32(-0.909743), f32(0.523083), f32(0.242386)],
			[f32(-0.747863), f32(0.22787), f32(-0.740794)],
			[f32(-0.678803), f32(-0.467344),
				f32(0.028562)],
			[f32(-0.11453), f32(0.564337), f32(0.910169)],
			[f32(0.11641), f32(-0.426091),
				f32(0.696344)],
			[f32(0.209231), f32(-0.02609), f32(-1.05619)],
			[f32(0.278291), f32(-0.721304),
				f32(-0.286836)],
			[f32(0.842564), f32(0.310377), f32(0.594771)],
			[f32(1.00444), f32(0.015163), f32(-0.38841)]]
		faces:    [[2, 6, 4], [6, 5, 8], [4, 7, 3], [2, 0, 1],
			[6, 2, 1, 5], [4, 6, 8, 7], [2, 4, 3, 0], [0, 3, 7, 8, 5, 1]]
	},
	&Polyhedron{
		name:     'j4'
		vertexes: [[f32(-0.600135), f32(0.398265), f32(-0.852158)],
			[f32(-0.585543), f32(-0.441941), f32(-0.840701)],
			[f32(-0.584691), f32(0.40999), f32(-0.011971)],
			[f32(-0.570099), f32(-0.430216),
				f32(-0.000514)],
			[f32(-0.18266), f32(1.00543), f32(-0.447988)],
			[f32(-0.147431), f32(-1.02301),
				f32(-0.420329)],
			[f32(0.0203), f32(0.428447), f32(0.571068)],
			[f32(0.034892), f32(-0.411759), f32(0.582525)],
			[f32(0.422331), f32(1.02389),
				f32(0.135052)],
			[f32(0.457559), f32(-1.00455), f32(0.162711)],
			[f32(0.860442), f32(0.442825),
				f32(0.555424)],
			[f32(0.875034), f32(-0.397381), f32(0.566881)]]
		faces:    [[3, 1, 5], [7, 9, 11], [6, 10, 8], [2, 4, 0],
			[2, 3, 7, 6], [3, 2, 0, 1], [7, 3, 5, 9], [6, 7, 11, 10],
			[2, 6, 8, 4], [4, 8, 10, 11, 9, 5, 1, 0]]
	},
	&Polyhedron{
		name:     'j5'
		vertexes: [[f32(-0.973114), f32(0.120196), f32(-0.57615)],
			[f32(-0.844191), f32(-0.563656), f32(-0.512814)],
			[f32(-0.711039), f32(0.75783), f32(-0.46202)],
			[f32(-0.594483), f32(0.244733),
				f32(-0.002202)],
			[f32(-0.46556), f32(-0.439119), f32(0.061133)],
			[f32(-0.373515), f32(-1.03252),
				f32(-0.296206)],
			[f32(-0.15807), f32(1.10569), f32(-0.21402)],
			[f32(-0.041514), f32(0.592595),
				f32(0.245798)],
			[f32(0.167087), f32(-0.513901), f32(0.348277)],
			[f32(0.259132), f32(-1.1073),
				f32(-0.009062)],
			[f32(0.429162), f32(0.123733), f32(0.462406)],
			[f32(0.474577), f32(1.03091), f32(0.073124)],
			[f32(0.812101), f32(-0.759438),
				f32(0.238938)],
			[f32(0.945253), f32(0.562048), f32(0.289732)],
			[f32(1.07418), f32(-0.121804),
				f32(0.353067)]]
		faces:    [[4, 1, 5], [8, 9, 12], [10, 14, 13], [7, 11, 6],
			[3, 2, 0], [4, 3, 0, 1], [8, 4, 5, 9], [10, 8, 12, 14],
			[7, 10, 13, 11], [3, 7, 6, 2], [3, 4, 8, 10, 7], [2, 6, 11, 13, 14, 12, 9, 5, 1, 0]]
	},
	&Polyhedron{
		name:     'j6'
		vertexes: [[f32(-0.905691), f32(-0.396105), f32(-0.539844)],
			[f32(-0.883472), f32(-0.258791), f32(0.103519)],
			[f32(-0.719735), f32(-0.859265),
				f32(-0.110695)],
			[f32(-0.703659), f32(0.13708), f32(-0.868724)],
			[f32(-0.667708), f32(0.359259),
				f32(0.17226)],
			[f32(-0.556577), f32(0.60392), f32(-0.428619)],
			[f32(-0.481752), f32(-0.103901),
				f32(0.60141)],
			[f32(-0.21682), f32(-1.07549), f32(0.254804)],
			[f32(-0.190808), f32(0.536633),
				f32(-0.971712)],
			[f32(-0.154857), f32(0.758811), f32(0.069272)],
			[f32(-0.069738), f32(-0.608646),
				f32(0.694909)],
			[f32(0.146026), f32(0.009404), f32(0.76365)],
			[f32(0.348059), f32(0.542589), f32(0.434771)],
			[f32(0.410958), f32(-0.962182),
				f32(0.417045)],
			[f32(0.436971), f32(0.649937), f32(-0.809472)],
			[f32(0.45919), f32(0.787251),
				f32(-0.166109)],
			[f32(0.760072), f32(0.037844), f32(0.52827)],
			[f32(0.923809), f32(-0.562629),
				f32(0.314056)],
			[f32(0.939886), f32(0.433715), f32(-0.443973)],
			[f32(1.12584), f32(-0.029444),
				f32(-0.014823)]]
		faces:    [[11, 16, 12], [16, 17, 19], [12, 15, 9], [15, 18, 14],
			[9, 5, 4], [5, 8, 3], [4, 1, 6], [1, 0, 2], [6, 10, 11],
			[10, 7, 13], [11, 12, 9, 4, 6], [11, 10, 13, 17, 16],
			[12, 16, 19, 18, 15], [9, 15, 14, 8, 5], [4, 5, 3, 0, 1],
			[6, 1, 2, 7, 10], [2, 0, 3, 8, 14, 18, 19, 17, 13, 7]]
	},
	&Polyhedron{
		name:     'j7'
		vertexes: [[f32(-0.793941), f32(-0.708614), f32(0.016702)],
			[f32(-0.451882), f32(0.284418), f32(0.56528)],
			[f32(-0.252303), f32(-0.348111),
				f32(-0.97361)],
			[f32(0.089756), f32(0.64492), f32(-0.425033)],
			[f32(0.340161), f32(-0.993103),
				f32(-0.175472)],
			[f32(0.385988), f32(1.12056), f32(0.619029)],
			[f32(0.68222), f32(-7.2e-05), f32(0.373105)]]
		faces:    [[0, 2, 4], [5, 3, 1], [5, 1, 6], [5, 6, 3],
			[3, 2, 0, 1], [1, 0, 4, 6], [6, 4, 2, 3]]
	},
	&Polyhedron{
		name:     'j8'
		vertexes: [[f32(-0.849167), f32(-0.427323), f32(0.457421)],
			[f32(-0.849167), f32(0.619869), f32(0.087182)],
			[f32(-0.478929), f32(-0.776386),
				f32(-0.529881)],
			[f32(-0.478929), f32(0.270805), f32(-0.900119)],
			[f32(0.198024), f32(-0.30391),
				f32(0.806484)],
			[f32(0.198024), f32(0.743282), f32(0.436246)],
			[f32(0.568263), f32(-0.652974),
				f32(-0.180817)],
			[f32(0.568263), f32(0.394218), f32(-0.551056)],
			[f32(1.12362), f32(0.13242), f32(0.37454)]]
		faces:    [[8, 7, 5], [8, 5, 4], [8, 4, 6], [8, 6, 7],
			[1, 3, 2, 0], [7, 3, 1, 5], [5, 1, 0, 4], [4, 0, 2, 6],
			[6, 2, 3, 7]]
	},
	&Polyhedron{
		name:     'j9'
		vertexes: [[f32(-0.980309), f32(-0.33878), f32(0.175213)],
			[f32(-0.719686), f32(0.629425), f32(0.02221)],
			[f32(-0.520232), f32(-0.599402),
				f32(-0.690328)],
			[f32(-0.299303), f32(-0.403757), f32(0.924054)],
			[f32(-0.25961), f32(0.368802),
				f32(-0.84333)],
			[f32(-0.03868), f32(0.564448), f32(0.771051)],
			[f32(0.243026), f32(0.902834),
				f32(-0.142672)],
			[f32(0.445117), f32(-0.825453), f32(-0.47642)],
			[f32(0.581659), f32(-0.704537),
				f32(0.521323)],
			[f32(0.705739), f32(0.142752), f32(-0.629422)],
			[f32(0.842281), f32(0.263667),
				f32(0.36832)]]
		faces:    [[6, 1, 5], [6, 5, 10], [6, 10, 9], [6, 9, 4],
			[6, 4, 1], [1, 0, 3, 5], [5, 3, 8, 10], [10, 8, 7, 9],
			[9, 7, 2, 4], [4, 2, 0, 1], [8, 3, 0, 2, 7]]
	},
	&Polyhedron{
		name:     'j10'
		vertexes: [[f32(-0.776892), f32(0.173498), f32(0.416855)],
			[f32(-0.68155), f32(0.270757), f32(-0.747914)],
			[f32(-0.646922), f32(-0.78715),
				f32(-0.243069)],
			[f32(0.020463), f32(0.897066), f32(-0.047806)],
			[f32(0.069435), f32(-0.599041),
				f32(0.666153)],
			[f32(0.15263), f32(0.505992), f32(1.04984)],
			[f32(0.480709), f32(0.236129), f32(-0.900199)],
			[f32(0.515337), f32(-0.821778),
				f32(-0.395353)],
			[f32(0.866791), f32(0.124527), f32(0.201492)]]
		faces:    [[4, 7, 8], [8, 7, 6], [8, 6, 3], [3, 6, 1],
			[3, 1, 0], [0, 1, 2], [0, 2, 4], [4, 2, 7], [4, 8, 5],
			[8, 3, 5], [3, 0, 5], [0, 4, 5], [1, 6, 7, 2]]
	},
	&Polyhedron{
		name:     'j11'
		vertexes: [[f32(-0.722759), f32(-0.425905), f32(0.628394)],
			[f32(-0.669286), f32(0.622275), f32(0.513309)],
			[f32(-0.502035), f32(-0.868253),
				f32(-0.304556)],
			[f32(-0.415513), f32(0.827739), f32(-0.490768)],
			[f32(-0.312146), f32(-0.093458),
				f32(-0.996236)],
			[f32(0.134982), f32(0.097675), f32(0.952322)],
			[f32(0.238349), f32(-0.823522),
				f32(0.446854)],
			[f32(0.324871), f32(0.872469), f32(0.260642)],
			[f32(0.492123), f32(-0.618058),
				f32(-0.557222)],
			[f32(0.545596), f32(0.430122), f32(-0.672308)],
			[f32(0.88582), f32(-0.021082),
				f32(0.21957)]]
		faces:    [[6, 2, 8], [8, 2, 4], [8, 4, 9], [9, 4, 3],
			[9, 3, 7], [7, 3, 1], [7, 1, 5], [5, 1, 0], [5, 0, 6],
			[6, 0, 2], [6, 8, 10], [8, 9, 10], [9, 7, 10], [7, 5, 10],
			[5, 6, 10], [1, 3, 4, 2, 0]]
	},
	&Polyhedron{
		name:     'j12'
		vertexes: [[f32(-0.610389), f32(0.243975), f32(0.531213)],
			[f32(-0.187812), f32(-0.48795), f32(-0.664016)],
			[f32(-0.187812), f32(0.9759),
				f32(-0.664016)],
			[f32(0.187812), f32(-0.9759), f32(0.664016)],
			[f32(0.798201), f32(0.243975), f32(0.132803)]]
		faces:    [[1, 3, 0], [3, 4, 0], [3, 1, 4], [0, 2, 1],
			[0, 4, 2], [2, 4, 1]]
	},
	&Polyhedron{
		name:     'j13'
		vertexes: [[f32(-1.02878), f32(0.392027), f32(-0.048786)],
			[f32(-0.640503), f32(-0.646161), f32(0.621837)],
			[f32(-0.125162), f32(-0.395663),
				f32(-0.540059)],
			[f32(0.004683), f32(0.888447), f32(-0.651988)],
			[f32(0.125161), f32(0.395663),
				f32(0.540059)],
			[f32(0.632925), f32(-0.791376), f32(0.433102)],
			[f32(1.03167), f32(0.157063),
				f32(-0.354165)]]
		faces:    [[3, 2, 0], [2, 1, 0], [2, 5, 1], [0, 4, 3],
			[0, 1, 4], [4, 1, 5], [2, 3, 6], [3, 4, 6], [5, 2, 6],
			[4, 5, 6]]
	},
	&Polyhedron{
		name:     'j14'
		vertexes: [[f32(-0.677756), f32(0.338878), f32(0.309352)],
			[f32(-0.446131), f32(1.33839), f32(0)], [f32(-0.338878), f32(-0.677755), f32(0.309352)],
			[f32(-0.169439), f32(0.508317), f32(-0.618703)],
			[f32(0.169439), f32(-0.508317),
				f32(-0.618703)],
			[f32(0.338878), f32(0.677756), f32(0.309352)], [f32(0.446131), f32(-1.33839), f32(0)],
			[f32(0.677755), f32(-0.338878), f32(0.309352)]]
		faces:    [[4, 7, 6], [5, 3, 1], [2, 4, 6], [3, 0, 1],
			[7, 2, 6], [0, 5, 1], [7, 4, 3, 5], [4, 2, 0, 3],
			[2, 7, 5, 0]]
	},
	&Polyhedron{
		name:     'j15'
		vertexes: [[f32(-0.669867), f32(0.334933), f32(-0.529576)],
			[f32(-0.669867), f32(0.334933), f32(0.529577)], [f32(-0.4043), f32(1.2129), f32(0)],
			[f32(-0.334933), f32(-0.669867), f32(-0.529576)],
			[f32(-0.334933), f32(-0.669867), f32(0.529577)],
			[f32(0.334933), f32(0.669867),
				f32(-0.529576)],
			[f32(0.334933), f32(0.669867), f32(0.529577)], [f32(0.4043), f32(-1.2129), f32(0)],
			[f32(0.669867), f32(-0.334933), f32(-0.529576)],
			[f32(0.669867), f32(-0.334933),
				f32(0.529577)]]
		faces:    [[8, 9, 7], [6, 5, 2], [3, 8, 7], [5, 0, 2],
			[4, 3, 7], [0, 1, 2], [9, 4, 7], [1, 6, 2], [9, 8, 5, 6],
			[8, 3, 0, 5], [3, 4, 1, 0], [4, 9, 6, 1]]
	},
	&Polyhedron{
		name:     'j16'
		vertexes: [[f32(-0.931836), f32(0.219976), f32(-0.264632)],
			[f32(-0.636706), f32(0.318353), f32(0.692816)],
			[f32(-0.613483), f32(-0.735083),
				f32(-0.264632)],
			[f32(-0.326545), f32(0.979634), f32(0)], [f32(-0.318353), f32(-0.636706), f32(0.692816)],
			[f32(-0.159176), f32(0.477529), f32(-0.856368)],
			[f32(0.159176), f32(-0.477529),
				f32(-0.856368)],
			[f32(0.318353), f32(0.636706), f32(0.692816)], [f32(0.326545), f32(-0.979634), f32(0)],
			[f32(0.613482), f32(0.735082), f32(-0.264632)],
			[f32(0.636706), f32(-0.318353),
				f32(0.692816)],
			[f32(0.931835), f32(-0.219977), f32(-0.264632)]]
		faces:    [[11, 10, 8], [7, 9, 3], [6, 11, 8], [9, 5, 3],
			[2, 6, 8], [5, 0, 3], [4, 2, 8], [0, 1, 3], [10, 4, 8],
			[1, 7, 3], [10, 11, 9, 7], [11, 6, 5, 9], [6, 2, 0, 5],
			[2, 4, 1, 0], [4, 10, 7, 1]]
	},
	&Polyhedron{
		name:     'j17'
		vertexes: [[f32(-0.777261), f32(0.485581), f32(0.103065)],
			[f32(-0.675344), f32(-0.565479), f32(-0.273294)],
			[f32(-0.379795), f32(-0.315718), f32(0.778861)],
			[f32(-0.221894), f32(0.282623),
				f32(-0.849372)],
			[f32(-0.034619), f32(1.23156), f32(-0.282624)],
			[f32(0.034619), f32(-1.23156),
				f32(0.282624)],
			[f32(0.196076), f32(0.635838), f32(0.638599)],
			[f32(0.405612), f32(-0.602744),
				f32(-0.568088)],
			[f32(0.701162), f32(-0.352983), f32(0.484067)],
			[f32(0.751443), f32(0.43288),
				f32(-0.313837)]]
		faces:    [[6, 8, 9], [9, 8, 7], [9, 7, 3], [3, 7, 1],
			[3, 1, 0], [0, 1, 2], [0, 2, 6], [6, 2, 8], [6, 9, 4],
			[9, 3, 4], [3, 0, 4], [0, 6, 4], [7, 8, 5], [1, 7, 5],
			[2, 1, 5], [8, 2, 5]]
	},
	&Polyhedron{
		name:     'j18'
		vertexes: [[f32(-0.836652), f32(0.050764), f32(0.288421)],
			[f32(-0.686658), f32(0.016522), f32(-0.560338)],
			[f32(-0.587106), f32(-0.771319),
				f32(0.365687)],
			[f32(-0.571616), f32(0.871513), f32(0.302147)],
			[f32(-0.437112), f32(-0.805561),
				f32(-0.483073)],
			[f32(-0.421621), f32(0.837272), f32(-0.546612)],
			[f32(-0.212729), f32(-0.16003),
				f32(0.84551)],
			[f32(0.052308), f32(0.660719), f32(0.859236)],
			[f32(0.08726), f32(-0.228514),
				f32(-0.852008)],
			[f32(0.186811), f32(-1.01636), f32(0.074016)],
			[f32(0.352296), f32(0.592236),
				f32(-0.838282)],
			[f32(0.561189), f32(-0.405066), f32(0.55384)],
			[f32(0.711183), f32(-0.439308),
				f32(-0.294919)],
			[f32(0.826226), f32(0.415684), f32(0.567566)],
			[f32(0.97622), f32(0.381442),
				f32(-0.281193)]]
		faces:    [[4, 9, 2], [9, 12, 11], [2, 6, 0], [4, 1, 8],
			[0, 3, 5, 1], [1, 5, 10, 8], [8, 10, 14, 12], [12, 14, 13, 11],
			[11, 13, 7, 6], [6, 7, 3, 0], [9, 4, 8, 12], [2, 9, 11, 6],
			[4, 2, 0, 1], [14, 10, 5, 3, 7, 13]]
	},
	&Polyhedron{
		name:     'j19'
		vertexes: [[f32(-0.889715), f32(0.115789), f32(-0.35951)],
			[f32(-0.792371), f32(-0.231368), f32(0.270291)],
			[f32(-0.791598), f32(0.494102),
				f32(0.251959)],
			[f32(-0.522446), f32(-0.406626), f32(-0.70424)],
			[f32(-0.521352), f32(0.619343),
				f32(-0.730164)],
			[f32(-0.425102), f32(-0.753782), f32(-0.074439)],
			[f32(-0.423235), f32(0.997655), f32(-0.118694)],
			[f32(-0.286344), f32(-0.218767),
				f32(0.790309)],
			[f32(-0.28557), f32(0.506702), f32(0.771978)],
			[f32(-0.154083), f32(0.096928),
				f32(-1.07489)],
			[f32(0.080926), f32(-0.741182), f32(0.44558)],
			[f32(0.082793), f32(1.01026), f32(0.401324)],
			[f32(0.095069), f32(-0.767118),
				f32(-0.580291)],
			[f32(0.331944), f32(0.146209), f32(0.895926)],
			[f32(0.463432), f32(-0.263565),
				f32(-0.950945)],
			[f32(0.601096), f32(-0.754518), f32(-0.060273)],
			[f32(0.699213), f32(-0.376205),
				f32(0.551197)],
			[f32(0.700307), f32(0.649763), f32(0.525272)],
			[f32(0.969459), f32(-0.250964),
				f32(-0.430927)],
			[f32(1.06758), f32(0.127349), f32(0.180543)]]
		faces:    [[10, 15, 16], [7, 13, 8], [1, 2, 0], [5, 3, 12],
			[2, 6, 4, 0], [0, 4, 9, 3], [3, 9, 14, 12], [12, 14, 18, 15],
			[15, 18, 19, 16], [16, 19, 17, 13], [13, 17, 11, 8],
			[8, 11, 6, 2], [5, 10, 7, 1], [10, 5, 12, 15], [7, 10, 16, 13],
			[1, 7, 8, 2], [5, 1, 0, 3], [18, 14, 9, 4, 6, 11, 17, 19]]
	},
	&Polyhedron{
		name:     'j20'
		vertexes: [[f32(-0.93465), f32(0.300459), f32(-0.271185)],
			[f32(-0.838689), f32(-0.260219), f32(-0.516017)],
			[f32(-0.711319), f32(0.717591), f32(0.128359)],
			[f32(-0.710334), f32(-0.156922),
				f32(0.080946)],
			[f32(-0.599799), f32(0.556003), f32(-0.725148)],
			[f32(-0.503838), f32(-0.004675),
				f32(-0.969981)],
			[f32(-0.487004), f32(0.26021), f32(0.48049)],
			[f32(-0.460089), f32(-0.750282),
				f32(-0.512622)],
			[f32(-0.376468), f32(0.973135), f32(-0.325605)],
			[f32(-0.331735), f32(-0.646985),
				f32(0.084342)],
			[f32(-0.254001), f32(0.831847), f32(0.530001)],
			[f32(-0.125239), f32(-0.494738),
				f32(-0.966586)],
			[f32(0.029622), f32(0.027949), f32(0.730817)],
			[f32(0.056536), f32(-0.982543),
				f32(-0.262295)],
			[f32(0.08085), f32(1.08739), f32(0.076037)],
			[f32(0.125583), f32(-0.532729), f32(0.485984)],
			[f32(0.262625), f32(0.599586),
				f32(0.780328)],
			[f32(0.391387), f32(-0.726999), f32(-0.716259)],
			[f32(0.513854), f32(-0.868287),
				f32(0.139347)],
			[f32(0.597475), f32(0.85513), f32(0.326364)],
			[f32(0.641224), f32(0.109523), f32(0.783723)],
			[f32(0.737185), f32(-0.451155),
				f32(0.538891)],
			[f32(0.848705), f32(-0.612742), f32(-0.314616)],
			[f32(0.976075), f32(0.365067),
				f32(0.32976)],
			[f32(1.07204), f32(-0.19561), f32(0.084927)]]
		faces:    [[15, 18, 21], [12, 20, 16], [6, 10, 2], [3, 0, 1],
			[9, 7, 13], [2, 8, 4, 0], [0, 4, 5, 1], [1, 5, 11, 7],
			[7, 11, 17, 13], [13, 17, 22, 18], [18, 22, 24, 21],
			[21, 24, 23, 20], [20, 23, 19, 16], [16, 19, 14, 10],
			[10, 14, 8, 2], [15, 9, 13, 18], [12, 15, 21, 20],
			[6, 12, 16, 10], [3, 6, 2, 0], [9, 3, 1, 7], [9, 15, 12, 6, 3],
			[22, 17, 11, 5, 4, 8, 14, 19, 23, 24]]
	},
	&Polyhedron{
		name:     'j21'
		vertexes: [[f32(-0.913903), f32(0.139054), f32(-0.10769)],
			[f32(-0.801323), f32(0.048332), f32(0.456301)],
			[f32(-0.780136), f32(-0.347362),
				f32(-0.398372)],
			[f32(-0.694081), f32(0.568652), f32(0.218063)],
			[f32(-0.672895), f32(0.172957),
				f32(-0.63661)],
			[f32(-0.597978), f32(-0.494154), f32(0.514184)],
			[f32(-0.584884), f32(-0.738707),
				f32(-0.014032)],
			[f32(-0.468218), f32(-0.603725), f32(-0.817867)],
			[f32(-0.378156), f32(-0.064556), f32(0.839937)],
			[f32(-0.360976), f32(-0.083405),
				f32(-1.05611)],
			[f32(-0.317215), f32(0.86806), f32(-0.109531)],
			[f32(-0.304122), f32(0.623508),
				f32(-0.637747)],
			[f32(-0.272966), f32(-0.995069), f32(-0.433527)],
			[f32(-0.204636), f32(0.777338), f32(0.45446)],
			[f32(-0.161718), f32(-0.851595),
				f32(0.369604)],
			[f32(-0.009384), f32(0.385994), f32(0.8388)],
			[f32(0.007796), f32(0.367145), f32(-1.05724)],
			[f32(0.1502), f32(-1.10796), f32(-0.049891)],
			[f32(0.185324), f32(0.832194), f32(-0.40135)],
			[f32(0.193961), f32(-0.156492),
				f32(0.896684)],
			[f32(0.327727), f32(-0.642909), f32(0.606002)],
			[f32(0.367482), f32(0.685403),
				f32(0.511206)],
			[f32(0.497242), f32(0.575832), f32(-0.820845)],
			[f32(0.60849), f32(0.719306),
				f32(-0.017714)],
			[f32(0.639645), f32(-0.899271), f32(0.186507)],
			[f32(0.6965), f32(-0.192358),
				f32(0.604864)],
			[f32(0.803742), f32(0.327961), f32(0.366626)],
			[f32(0.920408), f32(0.462943),
				f32(-0.437208)],
			[f32(1.00842), f32(-0.44872), f32(0.185369)],
			[f32(1.11566), f32(0.071599), f32(-0.052869)]]
		faces:    [[8, 19, 15], [19, 20, 25], [15, 21, 13], [21, 26, 23],
			[13, 10, 3], [10, 18, 11], [3, 0, 1], [0, 4, 2], [1, 5, 8],
			[5, 6, 14], [11, 16, 9, 4], [4, 9, 7, 2], [2, 7, 12, 6],
			[6, 12, 17, 14], [14, 17, 24, 20], [20, 24, 28, 25],
			[25, 28, 29, 26], [26, 29, 27, 23], [23, 27, 22, 18],
			[18, 22, 16, 11], [8, 15, 13, 3, 1], [8, 5, 14, 20, 19],
			[15, 19, 25, 26, 21], [13, 21, 23, 18, 10], [3, 10, 11, 4, 0],
			[1, 0, 2, 6, 5], [24, 17, 12, 7, 9, 16, 22, 27, 29, 28]]
	},
	&Polyhedron{
		name:     'j22'
		vertexes: [[f32(-0.846878), f32(0.066004), f32(0.311423)],
			[f32(-0.766106), f32(0.678635), f32(-0.329908)],
			[f32(-0.708152), f32(-0.186985),
				f32(-0.531132)],
			[f32(-0.64897), f32(-0.782761), f32(0.128183)],
			[f32(-0.452751), f32(0.845109),
				f32(0.48694)],
			[f32(-0.21247), f32(0.406919), f32(-0.972407)],
			[f32(-0.165405), f32(0.101357),
				f32(0.883692)],
			[f32(0.032503), f32(-0.747408), f32(0.700451)],
			[f32(0.112048), f32(-0.404621),
				f32(-0.801418)],
			[f32(0.17123), f32(-1.0004), f32(-0.142104)], [f32(0.41424), f32(0.739868), f32(0.66129)],
			[f32(0.654521), f32(0.301678), f32(-0.798058)],
			[f32(0.654794), f32(-0.116279),
				f32(0.613406)],
			[f32(0.793521), f32(-0.369268), f32(-0.229149)],
			[f32(0.967876), f32(0.468152),
				f32(0.018791)]]
		faces:    [[0, 1, 2], [2, 1, 5], [2, 5, 8], [8, 5, 11],
			[8, 11, 13], [13, 11, 14], [3, 9, 7], [9, 8, 13],
			[7, 12, 6], [3, 0, 2], [13, 14, 12], [12, 14, 10],
			[12, 10, 6], [6, 10, 4], [6, 4, 0], [0, 4, 1], [9, 3, 2, 8],
			[7, 9, 13, 12], [3, 7, 6, 0], [11, 5, 1, 4, 10, 14]]
	},
	&Polyhedron{
		name:     'j23'
		vertexes: [[f32(-0.96917), f32(0.321358), f32(-0.364138)],
			[f32(-0.902194), f32(0.146986), f32(0.353054)],
			[f32(-0.885918), f32(-0.386527),
				f32(-0.161101)],
			[f32(-0.700663), f32(0.819184), f32(0.114745)],
			[f32(-0.670588), f32(-0.166619),
				f32(-0.835289)],
			[f32(-0.389781), f32(0.533335), f32(0.723761)],
			[f32(-0.377102), f32(-0.207546),
				f32(0.737557)],
			[f32(-0.360826), f32(-0.741059), f32(0.223402)],
			[f32(-0.350486), f32(-0.754679),
				f32(-0.51752)],
			[f32(-0.022354), f32(1.03524), f32(0.320838)],
			[f32(0.020179), f32(-0.358897),
				f32(-1.02271)],
			[f32(0.351157), f32(0.546203), f32(0.733864)],
			[f32(0.363836), f32(-0.194678),
				f32(0.74766)],
			[f32(0.380112), f32(-0.728191), f32(0.233505)],
			[f32(0.390452), f32(-0.741811),
				f32(-0.507416)],
			[f32(0.668412), f32(0.842961), f32(0.133414)],
			[f32(0.698487), f32(-0.142842),
				f32(-0.816621)],
			[f32(0.886588), f32(0.178052), f32(0.377446)],
			[f32(0.902865), f32(-0.355461),
				f32(-0.136709)],
			[f32(0.966994), f32(0.354984), f32(-0.337737)]]
		faces:    [[1, 0, 2], [2, 0, 4], [2, 4, 8], [8, 4, 10],
			[8, 10, 14], [14, 10, 16], [14, 16, 18], [18, 16, 19],
			[13, 14, 18], [12, 17, 11], [6, 5, 1], [7, 2, 8],
			[18, 19, 17], [19, 15, 17], [17, 15, 11], [11, 15, 9],
			[11, 9, 5], [5, 9, 3], [5, 3, 1], [1, 3, 0], [7, 13, 12, 6],
			[13, 7, 8, 14], [12, 13, 18, 17], [6, 12, 11, 5],
			[7, 6, 1, 2], [10, 4, 0, 3, 9, 15, 19, 16]]
	},
	&Polyhedron{
		name:     'j24'
		vertexes: [[f32(-1.00794), f32(0.263193), f32(-0.317378)],
			[f32(-0.995648), f32(-0.249677), f32(0.04509)],
			[f32(-0.928425), f32(0.319026),
				f32(0.303212)],
			[f32(-0.878881), f32(-0.297121), f32(-0.570283)],
			[f32(-0.751014), f32(0.784617), f32(-0.079308)],
			[f32(-0.682946), f32(-0.746755),
				f32(-0.177844)],
			[f32(-0.534412), f32(-0.144902), f32(0.458433)],
			[f32(-0.506952), f32(0.74213),
				f32(0.497926)],
			[f32(-0.413141), f32(-0.682306), f32(-0.741423)],
			[f32(-0.221709), f32(-0.64198), f32(0.235499)],
			[f32(-0.206248), f32(1.06798),
				f32(0.052991)],
			[f32(-0.112939), f32(0.278202), f32(0.653148)],
			[f32(-0.109759), f32(-0.982341),
				f32(-0.280438)],
			[f32(0.107781), f32(0.858022), f32(0.55486)],
			[f32(0.211385), f32(-0.745233),
				f32(-0.765428)],
			[f32(0.393024), f32(-0.526088), f32(0.292433)],
			[f32(0.418278), f32(1.00506),
				f32(0.028986)],
			[f32(0.460247), f32(0.042616), f32(0.550554)],
			[f32(0.504974), f32(-0.866449),
				f32(-0.223504)],
			[f32(0.680968), f32(0.622436), f32(0.452266)],
			[f32(0.756151), f32(-0.461866),
				f32(-0.633128)],
			[f32(0.884017), f32(0.619872), f32(-0.142153)],
			[f32(0.926446), f32(-0.443346),
				f32(-0.028789)],
			[f32(0.99367), f32(0.125358), f32(0.229332)],
			[f32(1.01307), f32(0.059558), f32(-0.395059)]]
		faces:    [[1, 3, 5], [5, 3, 8], [5, 8, 12], [12, 8, 14],
			[12, 14, 18], [18, 14, 20], [18, 20, 22], [22, 20, 24],
			[22, 24, 23], [23, 24, 21], [15, 18, 22], [17, 23, 19],
			[11, 13, 7], [6, 2, 1], [9, 5, 12], [23, 21, 19],
			[19, 21, 16], [19, 16, 13], [13, 16, 10], [13, 10, 7],
			[7, 10, 4], [7, 4, 2], [2, 4, 0], [2, 0, 1], [1, 0, 3],
			[15, 9, 12, 18], [17, 15, 22, 23], [11, 17, 19, 13],
			[6, 11, 7, 2], [9, 6, 1, 5], [9, 15, 17, 11, 6], [20, 14, 8, 3, 0, 4, 10, 16, 21, 24]]
	},
	&Polyhedron{
		name:     'j25'
		vertexes: [[f32(-0.897802), f32(-0.193467), f32(-0.273331)],
			[f32(-0.877838), f32(-0.070089), f32(0.304735)],
			[f32(-0.73072), f32(-0.609618),
				f32(0.112262)],
			[f32(-0.716275), f32(0.285603), f32(-0.568831)],
			[f32(-0.703732), f32(-0.716856),
				f32(-0.46873)],
			[f32(-0.696138), f32(-0.246211), f32(-0.826802)],
			[f32(-0.683973), f32(0.485232), f32(0.366499)],
			[f32(-0.584121), f32(0.705062),
				f32(-0.173395)],
			[f32(-0.51689), f32(0.069081), f32(0.752092)],
			[f32(-0.378328), f32(-1.03778),
				f32(-0.09336)],
			[f32(-0.358446), f32(0.194389), f32(-1.0308)],
			[f32(-0.278847), f32(-0.803894),
				f32(0.440665)],
			[f32(-0.255475), f32(0.644603), f32(-0.661367)],
			[f32(-0.223173), f32(0.844232),
				f32(0.273963)],
			[f32(-0.146694), f32(-0.384435), f32(0.836102)],
			[f32(0.047172), f32(0.170886),
				f32(0.897866)],
			[f32(0.15578), f32(-1.08639), f32(0.15593)],
			[f32(0.180355), f32(0.436649), f32(-1.00282)],
			[f32(0.228699), f32(0.649956),
				f32(0.602366)],
			[f32(0.285215), f32(-0.70209), f32(0.586439)],
			[f32(0.308587), f32(0.746408),
				f32(-0.515593)],
			[f32(0.328551), f32(0.869786), f32(0.062473)],
			[f32(0.598896), f32(0.196439),
				f32(0.686376)],
			[f32(0.694582), f32(-0.844133), f32(0.183918)],
			[f32(0.714463), f32(0.388033),
				f32(-0.753526)],
			[f32(0.746014), f32(-0.343089), f32(0.493903)],
			[f32(0.760459), f32(0.552132),
				f32(-0.18719)],
			[f32(0.927542), f32(0.135981), f32(0.198403)],
			[f32(1.03227), f32(-0.403533),
				f32(-0.020084)],
			[f32(1.03987), f32(0.067112), f32(-0.378156)]]
		faces:    [[2, 9, 11], [11, 9, 16], [11, 16, 19], [19, 16, 23],
			[19, 23, 25], [25, 23, 28], [25, 28, 27], [27, 28, 29],
			[27, 29, 26], [26, 29, 24], [15, 22, 18], [22, 25, 27],
			[18, 21, 13], [21, 26, 20], [13, 7, 6], [7, 12, 3],
			[6, 1, 8], [1, 0, 2], [8, 14, 15], [14, 11, 19], [26, 24, 20],
			[20, 24, 17], [20, 17, 12], [12, 17, 10], [12, 10, 3],
			[3, 10, 5], [3, 5, 0], [0, 5, 4], [0, 4, 2], [2, 4, 9],
			[15, 18, 13, 6, 8], [15, 14, 19, 25, 22], [18, 22, 27, 26, 21],
			[13, 21, 20, 12, 7], [6, 7, 3, 0, 1], [8, 1, 2, 11, 14],
			[28, 23, 16, 9, 4, 5, 10, 17, 24, 29]]
	},
	&Polyhedron{
		name:     'j26'
		vertexes: [[f32(-0.57735), f32(0.57735), f32(0)], [f32(0.57735), f32(0.57735), f32(0)],
			[f32(0.57735), f32(-0.57735), f32(0)], [f32(-0.57735), f32(-0.57735), f32(0)],
			[f32(0), f32(0.57735), f32(1)], [f32(0), f32(-0.57735), f32(1)],
			[f32(-0.57735), f32(0), f32(-1)], [f32(0.57735), f32(0), f32(-1)]]
		faces:    [[1, 0, 4], [3, 2, 5], [3, 0, 6], [1, 2, 7],
			[3, 5, 4, 0], [1, 4, 5, 2], [1, 7, 6, 0], [3, 6, 7, 2]]
	},
	&Polyhedron{
		name:     'j27'
		vertexes: [[f32(-0.96936), f32(0.238651), f32(0.058198)],
			[f32(-0.683128), f32(-0.715413), f32(0.146701)],
			[f32(-0.623092), f32(-0.255511),
				f32(-0.739236)],
			[f32(-0.478567), f32(-0.06233), f32(0.875836)],
			[f32(-0.286232), f32(0.954064),
				f32(-0.088503)],
			[f32(0.060036), f32(0.459902), f32(-0.885938)],
			[f32(0.204561), f32(0.653083),
				f32(0.729135)],
			[f32(0.286232), f32(-0.954064), f32(0.088503)],
			[f32(0.346268), f32(-0.494162),
				f32(-0.797435)],
			[f32(0.490793), f32(-0.300981), f32(0.817638)],
			[f32(0.683128), f32(0.715413),
				f32(-0.146701)],
			[f32(0.96936), f32(-0.238651), f32(-0.058198)]]
		faces:    [[2, 5, 8], [5, 4, 10], [8, 11, 7], [2, 1, 0],
			[6, 3, 9], [3, 0, 1], [9, 7, 11], [6, 10, 4], [5, 2, 0, 4],
			[8, 5, 10, 11], [2, 8, 7, 1], [3, 6, 4, 0], [9, 3, 1, 7],
			[6, 9, 11, 10]]
	},
	&Polyhedron{
		name:     'j28'
		vertexes: [[f32(-1.0554), f32(0.383836), f32(-0.00011)],
			[f32(-1.01769), f32(-0.474869), f32(0.000238)],
			[f32(-0.474869), f32(1.01769),
				f32(-0.000394)],
			[f32(-0.448233), f32(0.410252), f32(-0.607929)],
			[f32(-0.448179), f32(0.410746),
				f32(0.607634)],
			[f32(-0.410526), f32(-0.448453), f32(-0.607581)],
			[f32(-0.410472), f32(-0.447959), f32(0.607981)],
			[f32(-0.383836), f32(-1.0554),
				f32(0.000446)],
			[f32(0.383836), f32(1.0554), f32(-0.000447)],
			[f32(0.410472), f32(0.447959),
				f32(-0.607982)],
			[f32(0.410526), f32(0.448453), f32(0.60758)],
			[f32(0.448179), f32(-0.410746),
				f32(-0.607635)],
			[f32(0.448233), f32(-0.410252), f32(0.607928)],
			[f32(0.474869), f32(-1.01769),
				f32(0.000392)],
			[f32(1.01769), f32(0.474869), f32(-0.000239)],
			[f32(1.0554), f32(-0.383836), f32(0.000109)]]
		faces:    [[3, 0, 2], [9, 8, 14], [11, 15, 13], [5, 7, 1],
			[6, 1, 7], [12, 13, 15], [10, 14, 8], [4, 2, 0], [5, 3, 9, 11],
			[3, 5, 1, 0], [9, 3, 2, 8], [11, 9, 14, 15], [5, 11, 13, 7],
			[4, 6, 12, 10], [6, 4, 0, 1], [12, 6, 7, 13], [10, 12, 15, 14],
			[4, 10, 8, 2]]
	},
	&Polyhedron{
		name:     'j29'
		vertexes: [[f32(-1.105), f32(-0.077473), f32(-0.184867)],
			[f32(-0.863019), f32(0.717824), f32(0.033637)],
			[f32(-0.699688), f32(-0.827387),
				f32(-0.295079)],
			[f32(-0.617244), f32(-0.39909), f32(0.445571)],
			[f32(-0.487757), f32(0.321617),
				f32(-0.630438)],
			[f32(-0.375262), f32(0.396206), f32(0.664075)],
			[f32(-0.115492), f32(1.09263),
				f32(0.232437)],
			[f32(-0.082444), f32(-0.428297), f32(-0.740649)],
			[f32(0.115493), f32(-1.09263), f32(-0.232437)],
			[f32(0.197937), f32(-0.664332),
				f32(0.508212)],
			[f32(0.25977), f32(0.696423), f32(-0.431638)],
			[f32(0.439918), f32(0.130964),
				f32(0.726716)],
			[f32(0.665082), f32(-0.053491), f32(-0.541849)],
			[f32(0.699688), f32(0.827387),
				f32(0.295079)],
			[f32(0.863019), f32(-0.717824), f32(-0.033637)],
			[f32(1.105), f32(0.077473), f32(0.184867)]]
		faces:    [[4, 0, 1], [10, 6, 13], [12, 15, 14], [7, 8, 2],
			[3, 0, 2], [9, 8, 14], [11, 15, 13], [5, 6, 1], [7, 4, 10, 12],
			[4, 7, 2, 0], [10, 4, 1, 6], [12, 10, 13, 15], [7, 12, 14, 8],
			[5, 3, 9, 11], [3, 5, 1, 0], [9, 3, 2, 8], [11, 9, 14, 15],
			[5, 11, 13, 6]]
	},
	&Polyhedron{
		name:     'j30'
		vertexes: [[f32(-1.19712), f32(-0.118752), f32(-0.001762)],
			[f32(-1.03824), f32(0.607337), f32(-0.020132)],
			[f32(-0.898745), f32(-0.799482),
				f32(0.017282)],
			[f32(-0.619431), f32(0.145275), f32(0.38469)],
			[f32(-0.61625), f32(0.124807),
				f32(-0.396793)],
			[f32(-0.482789), f32(1.10144), f32(-0.030813)],
			[f32(-0.321051), f32(-0.535454),
				f32(0.403734)],
			[f32(-0.317871), f32(-0.555923), f32(-0.37775)],
			[f32(-0.257075), f32(-1.17484),
				f32(0.029724)],
			[f32(-0.063976), f32(0.639383), f32(0.37401)],
			[f32(-0.060795), f32(0.618915),
				f32(-0.407474)],
			[f32(0.257076), f32(1.17484), f32(-0.029725)],
			[f32(0.418813), f32(-0.462061),
				f32(0.404823)],
			[f32(0.421993), f32(-0.48253), f32(-0.376661)],
			[f32(0.482789), f32(-1.10144),
				f32(0.030813)],
			[f32(0.577694), f32(0.264028), f32(0.386452)],
			[f32(0.580875), f32(0.24356),
				f32(-0.395032)],
			[f32(0.898745), f32(0.799482), f32(-0.017282)],
			[f32(1.03824), f32(-0.607337),
				f32(0.020132)],
			[f32(1.19712), f32(0.118752), f32(0.001761)]]
		faces:    [[4, 0, 1], [10, 5, 11], [16, 17, 19], [13, 18, 14],
			[7, 8, 2], [6, 2, 8], [12, 14, 18], [15, 19, 17],
			[9, 11, 5], [3, 1, 0], [4, 7, 2, 0], [10, 4, 1, 5],
			[16, 10, 11, 17], [13, 16, 19, 18], [7, 13, 14, 8],
			[6, 3, 0, 2], [12, 6, 8, 14], [15, 12, 18, 19], [9, 15, 17, 11],
			[3, 9, 5, 1], [7, 4, 10, 16, 13], [3, 6, 12, 15, 9]]
	},
	&Polyhedron{
		name:     'j31'
		vertexes: [[f32(-1.14213), f32(-0.353364), f32(-0.133745)],
			[f32(-1.13844), f32(0.385484), f32(-0.050817)],
			[f32(-0.70957), f32(-0.957238),
				f32(-0.165587)],
			[f32(-0.699897), f32(0.97709), f32(0.051522)],
			[f32(-0.598391), f32(0.052172),
				f32(-0.43817)],
			[f32(-0.543739), f32(-0.405536), f32(0.304426)],
			[f32(-0.540044), f32(0.333311),
				f32(0.387353)],
			[f32(-0.165831), f32(-0.551702), f32(-0.470012)],
			[f32(-0.159853), f32(0.643778), f32(-0.335832)],
			[f32(-0.005978), f32(-1.19548),
				f32(-0.13418)],
			[f32(0.005978), f32(1.19548), f32(0.134181)],
			[f32(0.159852), f32(-0.643778),
				f32(0.335832)],
			[f32(0.165831), f32(0.551702), f32(0.470012)],
			[f32(0.540044), f32(-0.333311),
				f32(-0.387353)],
			[f32(0.543739), f32(0.405536), f32(-0.304425)],
			[f32(0.598391), f32(-0.052172),
				f32(0.43817)],
			[f32(0.699896), f32(-0.97709), f32(-0.051521)],
			[f32(0.70957), f32(0.957238),
				f32(0.165587)],
			[f32(1.13844), f32(-0.385484), f32(0.050817)],
			[f32(1.14213), f32(0.353364), f32(0.133745)]]
		faces:    [[4, 0, 1], [8, 3, 10], [14, 17, 19], [13, 18, 16],
			[7, 9, 2], [5, 0, 2], [11, 9, 16], [15, 18, 19], [12, 17, 10],
			[6, 3, 1], [4, 7, 2, 0], [8, 4, 1, 3], [14, 8, 10, 17],
			[13, 14, 19, 18], [7, 13, 16, 9], [5, 6, 1, 0], [11, 5, 2, 9],
			[15, 11, 16, 18], [12, 15, 19, 17], [6, 12, 10, 3],
			[7, 4, 8, 14, 13], [6, 5, 11, 15, 12]]
	},
	&Polyhedron{
		name:     'j32'
		vertexes: [[f32(-1.08675), f32(0.270723), f32(-0.02221)],
			[f32(-0.951485), f32(0.016307), f32(0.590957)],
			[f32(-0.844123), f32(0.345447),
				f32(-0.65034)],
			[f32(-0.727726), f32(-0.227595), f32(-0.308179)],
			[f32(-0.678317), f32(0.606577), f32(0.401324)],
			[f32(-0.592457), f32(-0.482012),
				f32(0.304989)],
			[f32(-0.489983), f32(-0.320625), f32(0.954953)],
			[f32(-0.316268), f32(0.211936),
				f32(-1.05351)],
			[f32(-0.285732), f32(0.727482), f32(-0.61501)],
			[f32(-0.199871), f32(-0.361106),
				f32(-0.711346)],
			[f32(-0.183258), f32(0.888869), f32(0.034954)],
			[f32(-0.047989), f32(0.634452),
				f32(0.648121)],
			[f32(0.019), f32(-0.772761), f32(0.28078)], [f32(0.068408), f32(0.06141), f32(0.990283)],
			[f32(0.121473), f32(-0.611374), f32(0.930744)],
			[f32(0.261631), f32(-0.698037),
				f32(-0.34735)],
			[f32(0.295188), f32(-0.078813), f32(-1.07772)],
			[f32(0.344597), f32(0.755358),
				f32(-0.368213)],
			[f32(0.563468), f32(0.343703), f32(0.623912)],
			[f32(0.649328), f32(-0.744886),
				f32(0.527576)],
			[f32(0.703625), f32(0.25704), f32(-0.654181)],
			[f32(0.75669), f32(-0.415745),
				f32(-0.71372)],
			[f32(0.806099), f32(0.418427), f32(-0.004217)],
			[f32(0.891959), f32(-0.670162),
				f32(-0.100552)],
			[f32(0.922496), f32(-0.154616), f32(0.337944)]]
		faces:    [[3, 0, 2], [9, 7, 16], [15, 21, 23], [12, 19, 14],
			[5, 6, 1], [18, 24, 22], [24, 19, 23], [22, 20, 17],
			[20, 21, 16], [17, 8, 10], [8, 7, 2], [10, 4, 11],
			[4, 0, 1], [11, 13, 18], [13, 6, 14], [3, 5, 1, 0],
			[9, 3, 2, 7], [15, 9, 16, 21], [12, 15, 23, 19], [5, 12, 14, 6],
			[5, 3, 9, 15, 12], [18, 22, 17, 10, 11], [18, 13, 14, 19, 24],
			[22, 24, 23, 21, 20], [17, 20, 16, 7, 8], [10, 8, 2, 0, 4],
			[11, 4, 1, 6, 13]]
	},
	&Polyhedron{
		name:     'j33'
		vertexes: [[f32(-0.799512), f32(0.192706), f32(0.001565)],
			[f32(-0.776446), f32(0.593934), f32(0.546986)],
			[f32(-0.713384), f32(0.860598),
				f32(-0.072621)],
			[f32(-0.640335), f32(-0.34095), f32(0.387405)],
			[f32(-0.617268), f32(0.060277),
				f32(0.932827)],
			[f32(-0.538299), f32(0.090521), f32(-0.615141)],
			[f32(-0.452171), f32(0.758412),
				f32(-0.689327)],
			[f32(-0.296652), f32(-0.536533), f32(0.937522)],
			[f32(-0.280744), f32(-0.772953),
				f32(0.009162)],
			[f32(-0.217683), f32(-0.506289), f32(-0.610445)],
			[f32(-0.200278), f32(0.902051), f32(0.367837)],
			[f32(-0.09258), f32(0.326409),
				f32(-1.06757)],
			[f32(0.057277), f32(0.038576), f32(0.99214)],
			[f32(0.062939), f32(-0.968537),
				f32(0.559279)],
			[f32(0.222374), f32(0.736712), f32(-0.630014)],
			[f32(0.228036), f32(-0.270402),
				f32(-1.06287)],
			[f32(0.314991), f32(0.558821), f32(0.642957)],
			[f32(0.324152), f32(-1.07072),
				f32(-0.057426)],
			[f32(0.378052), f32(0.825485), f32(0.023349)],
			[f32(0.387214), f32(-0.804058),
				f32(-0.677033)],
			[f32(0.635607), f32(-0.037989), f32(0.647653)],
			[f32(0.639107), f32(-0.66042),
				f32(0.38013)],
			[f32(0.737643), f32(0.393482), f32(-0.354893)],
			[f32(0.741142), f32(-0.228948),
				f32(-0.622416)],
			[f32(0.89682), f32(-0.140175), f32(0.030947)]]
		faces:    [[5, 6, 11], [9, 15, 19], [8, 17, 13], [3, 7, 4],
			[0, 1, 2], [20, 21, 24], [21, 13, 17], [24, 23, 22],
			[23, 19, 15], [22, 14, 18], [14, 11, 6], [18, 10, 16],
			[10, 2, 1], [16, 12, 20], [12, 4, 7], [5, 0, 2, 6],
			[9, 5, 11, 15], [8, 9, 19, 17], [3, 8, 13, 7], [0, 3, 4, 1],
			[0, 5, 9, 8, 3], [20, 24, 22, 18, 16], [20, 12, 7, 13, 21],
			[24, 21, 17, 19, 23], [22, 23, 15, 11, 14], [18, 14, 6, 2, 10],
			[16, 10, 1, 4, 12]]
	},
	&Polyhedron{
		name:     'j34'
		vertexes: [[f32(-0.976027), f32(0.021192), f32(0.216616)],
			[f32(-0.8986), f32(-0.336852), f32(-0.281155)],
			[f32(-0.800821), f32(0.595002),
				f32(0.068255)],
			[f32(-0.778424), f32(-0.560713), f32(0.282236)],
			[f32(-0.680644), f32(0.371141),
				f32(0.631647)],
			[f32(-0.675542), f32(0.015675), f32(-0.737155)],
			[f32(-0.615111), f32(0.591592),
				f32(-0.521207)],
			[f32(-0.523949), f32(-0.823998), f32(-0.215648)],
			[f32(-0.360916), f32(-0.5704), f32(0.737823)],
			[f32(-0.319728), f32(0.941541),
				f32(-0.106177)],
			[f32(-0.300485), f32(0.005517), f32(0.953771)],
			[f32(-0.19445), f32(0.362214),
				f32(-0.911587)],
			[f32(-0.163033), f32(-0.253598), f32(-0.953472)],
			[f32(-0.125279), f32(0.579327), f32(0.80541)],
			[f32(-0.069344), f32(-0.772544),
				f32(-0.631163)],
			[f32(0.050833), f32(-0.996405), f32(-0.067772)],
			[f32(0.097779), f32(0.931854),
				f32(0.34941)],
			[f32(0.151593), f32(-0.839673), f32(0.521506)],
			[f32(0.194449), f32(-0.362214),
				f32(0.911587)],
			[f32(0.283489), f32(0.928444), f32(-0.240052)],
			[f32(0.360916), f32(0.5704),
				f32(-0.737823)],
			[f32(0.411749), f32(-0.426005), f32(-0.805595)],
			[f32(0.477939), f32(0.56623),
				f32(0.671534)],
			[f32(0.606198), f32(-0.788219), f32(0.105992)],
			[f32(0.675542), f32(-0.015675),
				f32(0.737155)],
			[f32(0.735567), f32(0.083254), f32(-0.672317)],
			[f32(0.778423), f32(0.560713),
				f32(-0.282236)],
			[f32(0.829257), f32(-0.435692), f32(-0.350008)],
			[f32(0.8986), f32(0.336852),
				f32(0.281155)],
			[f32(0.930017), f32(-0.27896),
				f32(0.23927)]]
		faces:    [[15, 7, 14], [7, 3, 1], [14, 12, 21], [12, 5, 11],
			[21, 25, 27], [25, 20, 26], [27, 29, 23], [29, 28, 24],
			[23, 17, 15], [17, 18, 8], [4, 10, 13], [10, 8, 18],
			[13, 22, 16], [22, 24, 28], [16, 19, 9], [19, 26, 20],
			[9, 6, 2], [6, 11, 5], [2, 0, 4], [0, 1, 3], [15, 14, 21, 27, 23],
			[15, 17, 8, 3, 7], [14, 7, 1, 5, 12], [21, 12, 11, 20, 25],
			[27, 25, 26, 28, 29], [23, 29, 24, 18, 17], [4, 13, 16, 9, 2],
			[4, 0, 3, 8, 10], [13, 10, 18, 24, 22], [16, 22, 28, 26, 19],
			[9, 19, 20, 11, 6], [2, 6, 5, 1, 0]]
	},
	&Polyhedron{
		name:     'j35'
		vertexes: [[f32(-0.903332), f32(-0.063468), f32(0.034076)],
			[f32(-0.833437), f32(0.28305), f32(0.763458)],
			[f32(-0.589483), f32(0.680853),
				f32(0.100738)],
			[f32(-0.561749), f32(-0.142046), f32(-0.696749)],
			[f32(-0.484641), f32(-0.705032), f32(0.29875)],
			[f32(-0.414746), f32(-0.358514),
				f32(1.02813)],
			[f32(-0.2479), f32(0.602275), f32(-0.630087)],
			[f32(-0.143058), f32(-0.78361),
				f32(-0.432074)],
			[f32(-0.100897), f32(0.385807), f32(1.09479)],
			[f32(0.065949), f32(0.076155), f32(-1.1608)],
			[f32(0.143058), f32(0.78361), f32(0.432075)],
			[f32(0.2479), f32(-0.602274), f32(0.630087)],
			[f32(0.484641), f32(-0.565409),
				f32(-0.896124)],
			[f32(0.484641), f32(0.705032), f32(-0.29875)],
			[f32(0.561749), f32(0.142046),
				f32(0.696749)],
			[f32(0.589483), f32(-0.680852), f32(-0.100737)],
			[f32(0.79849), f32(0.178912),
				f32(-0.829462)],
			[f32(0.903332), f32(0.063468), f32(-0.034075)]]
		faces:    [[9, 16, 12], [16, 13, 17], [12, 15, 7], [9, 3, 6],
			[8, 1, 5], [1, 2, 0], [5, 4, 11], [8, 14, 10], [16, 9, 6, 13],
			[12, 16, 17, 15], [9, 12, 7, 3], [1, 8, 10, 2], [5, 1, 0, 4],
			[8, 5, 11, 14], [7, 4, 0, 3], [3, 0, 2, 6], [6, 2, 10, 13],
			[13, 10, 14, 17], [17, 14, 11, 15], [15, 11, 4, 7]]
	},
	&Polyhedron{
		name:     'j36'
		vertexes: [[f32(-0.82124), f32(-0.196132), f32(-0.329082)],
			[f32(-0.725355), f32(-0.267867), f32(0.472553)],
			[f32(-0.627806), f32(0.589563),
				f32(-0.281911)],
			[f32(-0.577286), f32(0.20167), f32(-0.991803)],
			[f32(-0.531921), f32(0.517828),
				f32(0.519724)],
			[f32(-0.241376), f32(-0.749828), f32(-0.447988)],
			[f32(-0.196012), f32(-0.43367), f32(1.06354)],
			[f32(-0.145492), f32(-0.821562),
				f32(0.353647)],
			[f32(-0.002578), f32(0.352025), f32(1.11071)],
			[f32(0.002578), f32(-0.352025),
				f32(-1.11071)],
			[f32(0.145492), f32(0.821563), f32(-0.353646)],
			[f32(0.196012), f32(0.43367),
				f32(-1.06354)],
			[f32(0.241376), f32(0.749828), f32(0.447989)],
			[f32(0.531921), f32(-0.517828),
				f32(-0.519723)],
			[f32(0.577285), f32(-0.20167), f32(0.991804)],
			[f32(0.627806), f32(-0.589563),
				f32(0.281912)],
			[f32(0.725355), f32(0.267867), f32(-0.472551)],
			[f32(0.82124), f32(0.196133),
				f32(0.329083)]]
		faces:    [[3, 11, 9], [11, 10, 16], [9, 13, 5], [3, 0, 2],
			[14, 8, 6], [8, 12, 4], [6, 1, 7], [14, 15, 17], [11, 3, 2, 10],
			[9, 11, 16, 13], [3, 9, 5, 0], [8, 14, 17, 12], [6, 8, 4, 1],
			[14, 6, 7, 15], [5, 7, 1, 0], [0, 1, 4, 2], [2, 4, 12, 10],
			[10, 12, 17, 16], [16, 17, 15, 13], [13, 15, 7, 5]]
	},
	&Polyhedron{
		name:     'j37'
		vertexes: [[f32(-0.862856), f32(0.357407), f32(-0.357407)],
			[f32(-0.862856), f32(-0.357407), f32(-0.357407)],
			[f32(-0.357407), f32(0.862856), f32(-0.357407)],
			[f32(-0.357407), f32(0.357407),
				f32(-0.862856)],
			[f32(-0.357407), f32(-0.357407), f32(-0.862856)],
			[f32(-0.357407), f32(-0.862856), f32(-0.357407)],
			[f32(0.357407), f32(0.862856), f32(-0.357407)],
			[f32(0.357407), f32(0.357407),
				f32(-0.862856)],
			[f32(0.357407), f32(-0.357407), f32(-0.862856)],
			[f32(0.357407), f32(-0.862856),
				f32(-0.357407)],
			[f32(0.862856), f32(0.357407), f32(-0.357407)],
			[f32(0.862856), f32(-0.357407),
				f32(-0.357407)],
			[f32(0.862856), f32(0.357407), f32(0.357407)],
			[f32(0.862856), f32(-0.357407),
				f32(0.357407)],
			[f32(0.357407), f32(0.862856), f32(0.357407)], [f32(0.505449), f32(0), f32(0.862856)],
			[f32(0.357407), f32(-0.862856), f32(0.357407)], [f32(-0), f32(0.505449), f32(0.862856)],
			[f32(-0), f32(-0.505449), f32(0.862856)], [f32(-0.357407), f32(0.862856), f32(0.357407)],
			[f32(-0.505449), f32(0), f32(0.862856)], [f32(-0.357407), f32(-0.862856), f32(0.357407)],
			[f32(-0.862856), f32(0.357407), f32(0.357407)],
			[f32(-0.862856), f32(-0.357407),
				f32(0.357407)]]
		faces:    [[2, 3, 0], [4, 5, 1], [10, 7, 6], [11, 9, 8],
			[15, 13, 12], [19, 17, 14], [18, 21, 16], [22, 23, 20],
			[3, 4, 1, 0], [6, 7, 3, 2], [7, 8, 4, 3], [8, 9, 5, 4],
			[10, 11, 8, 7], [14, 17, 15, 12], [15, 18, 16, 13],
			[17, 20, 18, 15], [19, 22, 20, 17], [20, 23, 21, 18],
			[22, 19, 2, 0], [19, 14, 6, 2], [14, 12, 10, 6], [12, 13, 11, 10],
			[11, 13, 16, 9], [9, 16, 21, 5], [5, 21, 23, 1], [1, 23, 22, 0]]
	},
	&Polyhedron{
		name:     'j38'
		vertexes: [[f32(-1.04754), f32(-0.14473), f32(-0.164687)],
			[f32(-0.97266), f32(0.443085), f32(0.054945)],
			[f32(-0.794156), f32(0.029302),
				f32(-0.716846)],
			[f32(-0.77069), f32(-0.7105), f32(-0.215961)],
			[f32(-0.748241), f32(-0.047945),
				f32(0.383423)],
			[f32(-0.719275), f32(0.617116), f32(-0.497215)],
			[f32(-0.574648), f32(0.82842),
				f32(0.359043)],
			[f32(-0.517304), f32(-0.536469), f32(-0.76812)],
			[f32(-0.471389), f32(-0.613715),
				f32(0.332149)],
			[f32(-0.350229), f32(0.33739), f32(0.687521)],
			[f32(-0.321263), f32(1.00245),
				f32(-0.193117)],
			[f32(-0.247853), f32(-1.03812), f32(-0.079291)],
			[f32(-0.228431), f32(0.309073),
				f32(-0.749313)],
			[f32(-0.005532), f32(0.864089), f32(0.631452)],
			[f32(0.005532), f32(-0.864089),
				f32(-0.631452)],
			[f32(0.048421), f32(-0.256696), f32(-0.800587)],
			[f32(0.097726), f32(-0.578045),
				f32(0.604557)],
			[f32(0.169581), f32(0.694408), f32(-0.445215)],
			[f32(0.172608), f32(0.009769),
				f32(0.824189)],
			[f32(0.247853), f32(1.03812), f32(0.079291)],
			[f32(0.321263), f32(-1.00245), f32(0.193117)],
			[f32(0.517305), f32(0.536469), f32(0.76812)],
			[f32(0.574648), f32(-0.82842),
				f32(-0.359043)],
			[f32(0.617537), f32(-0.221027), f32(-0.528178)],
			[f32(0.692418), f32(0.366788),
				f32(-0.308546)],
			[f32(0.719275), f32(-0.617116), f32(0.497214)],
			[f32(0.77069), f32(0.7105), f32(0.215961)],
			[f32(0.794156), f32(-0.029301), f32(0.716846)],
			[f32(0.97266), f32(-0.443085),
				f32(-0.054945)],
			[f32(1.04754), f32(0.14473), f32(0.164687)]]
		faces:    [[17, 10, 19], [24, 26, 29], [23, 28, 22], [15, 14, 7],
			[12, 2, 5], [4, 1, 0], [8, 3, 11], [16, 20, 25], [18, 27, 21],
			[9, 13, 6], [17, 12, 5, 10], [24, 17, 19, 26], [23, 24, 29, 28],
			[15, 23, 22, 14], [12, 15, 7, 2], [4, 9, 6, 1], [8, 4, 0, 3],
			[16, 8, 11, 20], [18, 16, 25, 27], [9, 18, 21, 13],
			[22, 20, 11, 14], [14, 11, 3, 7], [7, 3, 0, 2], [2, 0, 1, 5],
			[5, 1, 6, 10], [10, 6, 13, 19], [19, 13, 21, 26],
			[26, 21, 27, 29], [29, 27, 25, 28], [28, 25, 20, 22],
			[12, 17, 24, 23, 15], [9, 4, 8, 16, 18]]
	},
	&Polyhedron{
		name:     'j39'
		vertexes: [[f32(-1.00686), f32(0.217224), f32(-0.290603)],
			[f32(-0.990318), f32(0.219795), f32(0.341133)],
			[f32(-0.944481), f32(-0.411647),
				f32(-0.289678)],
			[f32(-0.927935), f32(-0.409077), f32(0.342059)],
			[f32(-0.687819), f32(0.762632),
				f32(-0.301179)],
			[f32(-0.671273), f32(0.765203), f32(0.330558)],
			[f32(-0.551737), f32(-0.055664),
				f32(-0.63377)],
			[f32(-0.524499), f32(-0.883775), f32(-0.298756)],
			[f32(-0.507953), f32(-0.881203), f32(0.33298)],
			[f32(-0.446854), f32(0.274173),
				f32(0.659035)],
			[f32(-0.384471), f32(-0.354698), f32(0.65996)],
			[f32(-0.232692), f32(0.489744),
				f32(-0.644346)],
			[f32(-0.131755), f32(-0.527791), f32(-0.642848)],
			[f32(-0.10921), f32(1.01625), f32(-0.317365)],
			[f32(-0.092665), f32(1.01882),
				f32(0.314371)],
			[f32(0.092664), f32(-1.01882), f32(-0.314371)],
			[f32(0.10921), f32(-1.01625),
				f32(0.317365)],
			[f32(0.131755), f32(0.527791), f32(0.642848)],
			[f32(0.232692), f32(-0.489745),
				f32(0.644346)],
			[f32(0.384471), f32(0.354698), f32(-0.65996)],
			[f32(0.446854), f32(-0.274173),
				f32(-0.659035)],
			[f32(0.507953), f32(0.881203), f32(-0.33298)],
			[f32(0.524499), f32(0.883774),
				f32(0.298756)],
			[f32(0.551737), f32(0.055664), f32(0.63377)],
			[f32(0.671273), f32(-0.765203),
				f32(-0.330558)],
			[f32(0.687819), f32(-0.762632), f32(0.301179)],
			[f32(0.927935), f32(0.409076),
				f32(-0.342059)],
			[f32(0.944481), f32(0.411647), f32(0.289678)],
			[f32(0.990318), f32(-0.219795),
				f32(-0.341133)],
			[f32(1.00686), f32(-0.217224), f32(0.290603)]]
		faces:    [[11, 4, 13], [19, 21, 26], [20, 28, 24], [12, 15, 7],
			[6, 2, 0], [9, 5, 1], [10, 3, 8], [18, 16, 25], [23, 29, 27],
			[17, 22, 14], [11, 6, 0, 4], [19, 11, 13, 21], [20, 19, 26, 28],
			[12, 20, 24, 15], [6, 12, 7, 2], [9, 17, 14, 5], [10, 9, 1, 3],
			[18, 10, 8, 16], [23, 18, 25, 29], [17, 23, 27, 22],
			[24, 25, 16, 15], [15, 16, 8, 7], [7, 8, 3, 2], [2, 3, 1, 0],
			[0, 1, 5, 4], [4, 5, 14, 13], [13, 14, 22, 21], [21, 22, 27, 26],
			[26, 27, 29, 28], [28, 29, 25, 24], [6, 11, 19, 20, 12],
			[17, 9, 10, 18, 23]]
	},
	&Polyhedron{
		name:     'j40'
		vertexes: [[f32(-1.05518), f32(-0.061289), f32(-0.047893)],
			[f32(-0.934164), f32(0.280612), f32(0.409939)],
			[f32(-0.859454), f32(-0.241561),
				f32(-0.56784)],
			[f32(-0.777777), f32(-0.505581), f32(0.210572)],
			[f32(-0.776073), f32(0.311702),
				f32(-0.400212)],
			[f32(-0.656761), f32(-0.163679), f32(0.668404)],
			[f32(-0.655057), f32(0.653604),
				f32(0.05762)],
			[f32(-0.582051), f32(-0.685853), f32(-0.309375)],
			[f32(-0.542629), f32(0.653549), f32(0.63078)],
			[f32(-0.421745), f32(-0.191346),
				f32(-0.9513)],
			[f32(-0.400139), f32(-0.685942), f32(0.618017)],
			[f32(-0.338365), f32(0.361918),
				f32(-0.783672)],
			[f32(-0.265226), f32(0.209257), f32(0.889245)],
			[f32(-0.144342), f32(-0.635637),
				f32(-0.692835)],
			[f32(-0.142556), f32(0.915126), f32(-0.042884)],
			[f32(-0.083446), f32(-0.977628),
				f32(-0.223275)],
			[f32(-0.030129), f32(0.915071), f32(0.530275)],
			[f32(0.028982), f32(-0.977682),
				f32(0.349884)],
			[f32(0.05317), f32(0.734854), f32(-0.562831)],
			[f32(0.090755), f32(0.070177),
				f32(-1.05181)],
			[f32(0.149998), f32(-0.635781), f32(0.807716)],
			[f32(0.233378), f32(-0.082518),
				f32(0.975345)],
			[f32(0.247274), f32(0.47078), f32(0.788741)],
			[f32(0.368158), f32(-0.374115),
				f32(-0.793339)],
			[f32(0.40758), f32(0.965287), f32(0.146815)],
			[f32(0.46669), f32(-0.927467),
				f32(-0.033576)],
			[f32(0.48229), f32(0.443114), f32(-0.830964)],
			[f32(0.603306), f32(0.785015),
				f32(-0.373132)],
			[f32(0.662498), f32(-0.374258), f32(0.707212)],
			[f32(0.684983), f32(0.520995),
				f32(0.405281)],
			[f32(0.745797), f32(-0.554475), f32(-0.385895)],
			[f32(0.759693), f32(-0.001178),
				f32(-0.572498)],
			[f32(0.858225), f32(-0.55453), f32(0.187265)],
			[f32(0.880709), f32(0.340724),
				f32(-0.114666)],
			[f32(0.941605), f32(-0.001267), f32(0.354893)]]
		faces:    [[6, 1, 8], [14, 16, 24], [18, 27, 26], [11, 19, 9],
			[4, 2, 0], [20, 10, 17], [10, 5, 3], [17, 15, 25],
			[15, 7, 13], [25, 30, 32], [30, 23, 31], [32, 34, 28],
			[34, 33, 29], [28, 21, 20], [21, 22, 12], [6, 4, 0, 1],
			[14, 6, 8, 16], [18, 14, 24, 27], [11, 18, 26, 19],
			[4, 11, 9, 2], [26, 31, 23, 19], [19, 23, 13, 9],
			[9, 13, 7, 2], [2, 7, 3, 0], [0, 3, 5, 1], [1, 5, 12, 8],
			[8, 12, 22, 16], [16, 22, 29, 24], [24, 29, 33, 27],
			[27, 33, 31, 26], [4, 6, 14, 18, 11], [20, 17, 25, 32, 28],
			[20, 21, 12, 5, 10], [17, 10, 3, 7, 15], [25, 15, 13, 23, 30],
			[32, 30, 31, 33, 34], [28, 34, 29, 22, 21]]
	},
	&Polyhedron{
		name:     'j41'
		vertexes: [[f32(-1.04503), f32(0.161365), f32(0.036367)],
			[f32(-0.919366), f32(0.043922), f32(-0.521815)],
			[f32(-0.855707), f32(-0.369212),
				f32(0.190625)],
			[f32(-0.830432), f32(0.382234), f32(0.532668)],
			[f32(-0.73004), f32(-0.486655),
				f32(-0.367556)],
			[f32(-0.711442), f32(0.52894), f32(-0.271461)],
			[f32(-0.641106), f32(-0.148342),
				f32(0.686927)],
			[f32(-0.544409), f32(-0.844483), f32(0.055116)],
			[f32(-0.501432), f32(0.074765),
				f32(-0.928671)],
			[f32(-0.496841), f32(0.749809), f32(0.224841)],
			[f32(-0.357534), f32(0.622166),
				f32(0.777518)],
			[f32(-0.312106), f32(-0.455811), f32(-0.774412)],
			[f32(-0.293508), f32(0.559783), f32(-0.678317)],
			[f32(-0.197177), f32(-0.487108),
				f32(0.858148)],
			[f32(-0.168208), f32(0.09159), f32(0.931777)],
			[f32(-0.137415), f32(-0.917347),
				f32(0.467667)],
			[f32(-0.011748), f32(-1.03479), f32(-0.090514)],
			[f32(0.049132), f32(0.242114),
				f32(-1.0288)],
			[f32(0.053724), f32(0.917158), f32(0.124716)],
			[f32(0.131823), f32(-0.794577),
				f32(-0.603191)],
			[f32(0.17939), f32(0.799715), f32(-0.433466)],
			[f32(0.193031), f32(0.789515),
				f32(0.677394)],
			[f32(0.238459), f32(-0.288463), f32(-0.874537)],
			[f32(0.335483), f32(-0.677415),
				f32(0.712518)],
			[f32(0.382357), f32(0.258938), f32(0.831652)],
			[f32(0.522031), f32(0.482046),
				f32(-0.783946)],
			[f32(0.538816), f32(-0.867441), f32(-0.190639)],
			[f32(0.610965), f32(0.820358),
				f32(0.270538)],
			[f32(0.693655), f32(-0.216333), f32(0.696143)],
			[f32(0.711357), f32(-0.048531),
				f32(-0.629687)],
			[f32(0.736632), f32(0.702915), f32(-0.287644)],
			[f32(0.753417), f32(-0.646572),
				f32(0.305662)],
			[f32(0.800291), f32(0.289782), f32(0.424796)],
			[f32(0.896988), f32(-0.406359),
				f32(-0.207015)],
			[f32(0.925958), f32(0.172339), f32(-0.133386)]]
		faces:    [[9, 3, 10], [18, 21, 27], [20, 30, 25], [12, 17, 8],
			[5, 1, 0], [15, 7, 16], [7, 2, 4], [16, 19, 26], [19, 11, 22],
			[26, 33, 31], [33, 29, 34], [31, 28, 23], [28, 32, 24],
			[23, 13, 15], [13, 14, 6], [9, 5, 0, 3], [18, 9, 10, 21],
			[20, 18, 27, 30], [12, 20, 25, 17], [5, 12, 8, 1],
			[25, 29, 22, 17], [17, 22, 11, 8], [8, 11, 4, 1],
			[1, 4, 2, 0], [0, 2, 6, 3], [3, 6, 14, 10], [10, 14, 24, 21],
			[21, 24, 32, 27], [27, 32, 34, 30], [30, 34, 29, 25],
			[5, 9, 18, 20, 12], [15, 16, 26, 31, 23], [15, 13, 6, 2, 7],
			[16, 7, 4, 11, 19], [26, 19, 22, 29, 33], [31, 33, 34, 32, 28],
			[23, 28, 24, 14, 13]]
	},
	&Polyhedron{
		name:     'j42'
		vertexes: [[f32(-1.09423), f32(0.091579), f32(-0.183298)],
			[f32(-0.983491), f32(-0.29488), f32(0.177777)],
			[f32(-0.97462), f32(-0.408146),
				f32(-0.350504)],
			[f32(-0.882171), f32(0.554599), f32(-0.002654)],
			[f32(-0.873301), f32(0.441333),
				f32(-0.530935)],
			[f32(-0.702994), f32(-0.070704), f32(0.581578)],
			[f32(-0.679771), f32(-0.367238),
				f32(-0.801479)],
			[f32(-0.640375), f32(0.454303), f32(0.470066)],
			[f32(-0.617152), f32(0.157769),
				f32(-0.912991)],
			[f32(-0.583386), f32(-0.570429), f32(0.414373)],
			[f32(-0.569033), f32(-0.753697),
				f32(-0.440404)],
			[f32(-0.419447), f32(0.804058), f32(0.122429)],
			[f32(-0.405095), f32(0.620789),
				f32(-0.732347)],
			[f32(-0.327237), f32(-0.853993), f32(0.032316)],
			[f32(-0.251159), f32(-0.061675),
				f32(0.877809)],
			[f32(-0.211565), f32(-0.187782), f32(-1.00289)],
			[f32(-0.18854), f32(0.463332),
				f32(0.766296)],
			[f32(-0.131551), f32(-0.5614), f32(0.710603)],
			[f32(-0.124598), f32(0.844965),
				f32(-0.328546)],
			[f32(-0.032387), f32(-0.813085), f32(-0.41866)],
			[f32(0.032387), f32(0.813086),
				f32(0.418659)],
			[f32(0.124598), f32(-0.844964), f32(0.328546)],
			[f32(0.131551), f32(0.561401),
				f32(-0.710603)],
			[f32(0.18854), f32(-0.463331), f32(-0.766296)],
			[f32(0.237051), f32(-0.270491),
				f32(0.977985)],
			[f32(0.251159), f32(0.061676), f32(-0.877809)],
			[f32(0.327237), f32(0.853994),
				f32(-0.032316)],
			[f32(0.33837), f32(0.578988), f32(0.797554)],
			[f32(0.419448), f32(-0.804057),
				f32(-0.122429)],
			[f32(0.583386), f32(0.570429), f32(-0.414373)],
			[f32(0.601401), f32(0.125461),
				f32(0.928384)],
			[f32(0.640375), f32(-0.454302), f32(-0.470066)],
			[f32(0.651509), f32(-0.729308),
				f32(0.359803)],
			[f32(0.702994), f32(0.070705), f32(-0.581579)],
			[f32(0.721009), f32(-0.374264),
				f32(0.761179)],
			[f32(0.815447), f32(0.645178), f32(0.06786)],
			[f32(0.822328), f32(0.475215), f32(0.580748)],
			[f32(1.00898), f32(-0.163393),
				f32(-0.202684)],
			[f32(1.01586), f32(-0.333356), f32(0.310203)],
			[f32(1.07848), f32(0.191651), f32(0.198691)]]
		faces:    [[0, 3, 4], [3, 7, 11], [4, 12, 8], [12, 18, 22],
			[8, 15, 6], [15, 25, 23], [6, 10, 2], [10, 19, 13],
			[2, 1, 0], [1, 9, 5], [30, 24, 34], [24, 14, 17],
			[34, 32, 38], [32, 21, 28], [38, 37, 39], [37, 31, 33],
			[39, 35, 36], [35, 29, 26], [36, 27, 30], [27, 20, 16],
			[23, 31, 28, 19], [19, 28, 21, 13], [13, 21, 17, 9],
			[9, 17, 14, 5], [5, 14, 16, 7], [7, 16, 20, 11], [11, 20, 26, 18],
			[18, 26, 29, 22], [22, 29, 33, 25], [25, 33, 31, 23],
			[0, 4, 8, 6, 2], [0, 1, 5, 7, 3], [4, 3, 11, 18, 12],
			[8, 12, 22, 25, 15], [6, 15, 23, 19, 10], [2, 10, 13, 9, 1],
			[30, 34, 38, 39, 36], [30, 27, 16, 14, 24], [34, 24, 17, 21, 32],
			[38, 32, 28, 31, 37], [39, 37, 33, 29, 35], [36, 35, 26, 20, 27]]
	},
	&Polyhedron{
		name:     'j43'
		vertexes: [[f32(-1.09992), f32(-0.170755), f32(-0.018241)],
			[f32(-1.01574), f32(0.184543), f32(-0.41657)],
			[f32(-0.979069), f32(0.342745),
				f32(0.098809)],
			[f32(-0.891012), f32(-0.645186), f32(-0.17075)],
			[f32(-0.854337), f32(-0.486985),
				f32(0.344629)],
			[f32(-0.754806), f32(-0.070303), f32(-0.81526)],
			[f32(-0.677717), f32(-0.583103),
				f32(-0.663335)],
			[f32(-0.65879), f32(0.343875), f32(0.53402)],
			[f32(-0.633951), f32(0.443197),
				f32(-0.698209)],
			[f32(-0.581702), f32(-0.168926), f32(0.685945)],
			[f32(-0.57461), f32(0.699173),
				f32(0.135692)],
			[f32(-0.43213), f32(-0.899333), f32(-0.300465)],
			[f32(-0.37279), f32(-0.643357),
				f32(0.533436)],
			[f32(-0.361315), f32(0.761256), f32(-0.356893)],
			[f32(-0.295924), f32(-0.324449),
				f32(-0.944974)],
			[f32(-0.185624), f32(0.480819), f32(0.756166)],
			[f32(-0.111851), f32(-0.898203),
				f32(0.134746)],
			[f32(-0.108536), f32(-0.031982), f32(0.908091)],
			[f32(-0.101444), f32(0.836117),
				f32(0.357838)],
			[f32(-0.100377), f32(0.50641), f32(-0.755583)],
			[f32(0.100376), f32(-0.506413),
				f32(0.755582)],
			[f32(0.101443), f32(-0.83612), f32(-0.357838)],
			[f32(0.108535), f32(0.031979),
				f32(-0.908092)],
			[f32(0.111851), f32(0.8982), f32(-0.134747)],
			[f32(0.185623), f32(-0.480822),
				f32(-0.756167)],
			[f32(0.295923), f32(0.324447), f32(0.944974)],
			[f32(0.361314), f32(-0.761258),
				f32(0.356892)],
			[f32(0.372789), f32(0.643354), f32(-0.533437)],
			[f32(0.43213), f32(0.899331),
				f32(0.300464)],
			[f32(0.574609), f32(-0.699176), f32(-0.135692)],
			[f32(0.581701), f32(0.168923),
				f32(-0.685946)],
			[f32(0.63395), f32(-0.443199), f32(0.698208)],
			[f32(0.658789), f32(-0.343878),
				f32(-0.534021)],
			[f32(0.677716), f32(0.583101), f32(0.663334)],
			[f32(0.754804), f32(0.0703), f32(0.815259)],
			[f32(0.854336), f32(0.486982), f32(-0.344629)],
			[f32(0.891011), f32(0.645184),
				f32(0.17075)],
			[f32(0.979068), f32(-0.342747), f32(-0.09881)],
			[f32(1.01574), f32(-0.184545),
				f32(0.416569)],
			[f32(1.09992), f32(0.170753), f32(0.018241)]]
		faces:    [[0, 2, 1], [2, 7, 10], [1, 8, 5], [8, 13, 19],
			[5, 14, 6], [14, 22, 24], [6, 11, 3], [11, 21, 16],
			[3, 4, 0], [4, 12, 9], [33, 25, 34], [25, 15, 17],
			[34, 31, 38], [31, 20, 26], [38, 37, 39], [37, 29, 32],
			[39, 35, 36], [35, 30, 27], [36, 28, 33], [28, 23, 18],
			[24, 32, 29, 21], [21, 29, 26, 16], [16, 26, 20, 12],
			[12, 20, 17, 9], [9, 17, 15, 7], [7, 15, 18, 10],
			[10, 18, 23, 13], [13, 23, 27, 19], [19, 27, 30, 22],
			[22, 30, 32, 24], [0, 1, 5, 6, 3], [0, 4, 9, 7, 2],
			[1, 2, 10, 13, 8], [5, 8, 19, 22, 14], [6, 14, 24, 21, 11],
			[3, 11, 16, 12, 4], [33, 34, 38, 39, 36], [33, 28, 18, 15, 25],
			[34, 25, 17, 20, 31], [38, 31, 26, 29, 37], [39, 37, 32, 30, 35],
			[36, 35, 27, 23, 28]]
	},
	&Polyhedron{
		name:     'j44'
		vertexes: [[f32(-0.789003), f32(0.385273), f32(-0.254111)],
			[f32(-0.772339), f32(-0.452189), f32(-0.185879)],
			[f32(-0.761383), f32(0.026005), f32(0.505125)],
			[f32(-0.611639), f32(-0.798949),
				f32(0.562592)],
			[f32(-0.381598), f32(-0.074991), f32(-0.82722)],
			[f32(-0.362623), f32(0.753266),
				f32(0.369634)],
			[f32(-0.289802), f32(0.760316), f32(-0.816621)],
			[f32(-0.055737), f32(-0.771195),
				f32(-0.487529)],
			[f32(-0.033826), f32(0.185193), f32(0.894479)],
			[f32(0.104963), f32(-1.11796),
				f32(0.260942)],
			[f32(0.115918), f32(-0.639761), f32(0.951946)],
			[f32(0.136578), f32(1.12831),
				f32(-0.192876)],
			[f32(0.452187), f32(-0.167262), f32(-0.776585)],
			[f32(0.471162), f32(0.660994),
				f32(0.420269)],
			[f32(0.543983), f32(0.668044), f32(-0.765985)],
			[f32(0.67182), f32(-0.612007),
				f32(-0.098176)],
			[f32(0.682775), f32(-0.133813), f32(0.592828)],
			[f32(0.878567), f32(0.200731),
				f32(-0.15284)]]
		faces:    [[11, 14, 6], [14, 17, 12], [6, 4, 0], [11, 5, 13],
			[9, 10, 3], [10, 16, 8], [3, 2, 1], [9, 7, 15], [4, 1, 0],
			[0, 1, 2], [0, 2, 5], [5, 2, 8], [5, 8, 13], [13, 8, 16],
			[13, 16, 17], [17, 16, 15], [17, 15, 12], [12, 15, 7],
			[12, 7, 4], [4, 7, 1], [14, 11, 13, 17], [6, 14, 12, 4],
			[11, 6, 0, 5], [10, 9, 15, 16], [3, 10, 8, 2], [9, 3, 1, 7]]
	},
	&Polyhedron{
		name:     'j45'
		vertexes: [[f32(-0.984615), f32(-0.215433), f32(0.042813)],
			[f32(-0.835086), f32(0.417027), f32(0.382665)],
			[f32(-0.776626), f32(0.078669),
				f32(-0.596021)],
			[f32(-0.681291), f32(-0.220722), f32(0.710519)],
			[f32(-0.642753), f32(-0.628915),
				f32(-0.457214)],
			[f32(-0.627097), f32(0.71113), f32(-0.256169)],
			[f32(-0.577202), f32(-0.786781),
				f32(0.255979)],
			[f32(-0.300907), f32(0.381853), f32(0.883943)],
			[f32(-0.281757), f32(0.897979),
				f32(0.36326)],
			[f32(-0.143631), f32(0.126378), f32(-0.963315)],
			[f32(-0.068623), f32(-0.621064),
				f32(0.757726)],
			[f32(-0.049613), f32(-0.984736), f32(-0.213412)],
			[f32(-0.009758), f32(-0.581206), f32(-0.824509)],
			[f32(0.005899), f32(0.758839), f32(-0.623463)],
			[f32(0.311761), f32(-0.018489),
				f32(0.931151)],
			[f32(0.341127), f32(0.667962), f32(0.674663)],
			[f32(0.351238), f32(0.945688),
				f32(-0.004035)],
			[f32(0.458966), f32(-0.819019), f32(0.288335)],
			[f32(0.54357), f32(-0.100253),
				f32(-0.843914)],
			[f32(0.592421), f32(-0.698626), f32(-0.422693)],
			[f32(0.6931), f32(0.532207),
				f32(-0.504062)],
			[f32(0.83935), f32(-0.216444), f32(0.461759)],
			[f32(0.868716), f32(0.470008),
				f32(0.205272)],
			[f32(0.972805), f32(-0.096052), f32(-0.249268)]]
		faces:    [[13, 16, 20], [9, 18, 12], [2, 4, 0], [5, 1, 8],
			[14, 15, 7], [10, 3, 6], [17, 11, 19], [21, 23, 22],
			[12, 11, 4], [4, 11, 6], [4, 6, 0], [0, 6, 3], [0, 3, 1],
			[1, 3, 7], [1, 7, 8], [8, 7, 15], [8, 15, 16], [16, 15, 22],
			[16, 22, 20], [20, 22, 23], [20, 23, 18], [18, 23, 19],
			[18, 19, 12], [12, 19, 11], [5, 13, 9, 2], [13, 5, 8, 16],
			[9, 13, 20, 18], [2, 9, 12, 4], [5, 2, 0, 1], [21, 14, 10, 17],
			[14, 21, 22, 15], [10, 14, 7, 3], [17, 10, 6, 11],
			[21, 17, 19, 23]]
	},
	&Polyhedron{
		name:     'j46'
		vertexes: [[f32(-0.962816), f32(0.187793), f32(0.445444)],
			[f32(-0.942301), f32(-0.435696), f32(0.287991)],
			[f32(-0.736715), f32(0.34226),
				f32(-0.136766)],
			[f32(-0.7162), f32(-0.281228), f32(-0.294218)],
			[f32(-0.680334), f32(0.758077),
				f32(0.35095)],
			[f32(-0.653736), f32(-0.229833), f32(0.824928)],
			[f32(-0.626624), f32(-0.874236),
				f32(-0.061265)],
			[f32(-0.516012), f32(0.397771), f32(0.858028)],
			[f32(-0.47699), f32(-0.788175),
				f32(0.558536)],
			[f32(-0.259134), f32(0.641512), f32(-0.447112)],
			[f32(-0.22594), f32(-0.367313),
				f32(-0.701875)],
			[f32(-0.202753), f32(1.05733), f32(0.040605)],
			[f32(-0.136364), f32(-0.960322),
				f32(-0.468922)],
			[f32(-0.116423), f32(0.854913), f32(0.645191)],
			[f32(-0.053283), f32(-1.06399),
				f32(0.160603)],
			[f32(-0.029965), f32(-0.362198), f32(0.739264)],
			[f32(0.056543), f32(0.202971),
				f32(-0.796368)],
			[f32(0.107759), f32(0.265405), f32(0.772363)],
			[f32(0.287508), f32(0.971244),
				f32(-0.367052)],
			[f32(0.341218), f32(-0.66107), f32(-0.779268)],
			[f32(0.392401), f32(0.966981),
				f32(0.267715)],
			[f32(0.393741), f32(-0.638011), f32(0.341331)],
			[f32(0.455541), f32(-0.951919),
				f32(-0.216873)],
			[f32(0.603185), f32(0.532703), f32(-0.716309)],
			[f32(0.616584), f32(0.377473),
				f32(0.394887)],
			[f32(0.6237), f32(-0.090786), f32(-0.873761)],
			[f32(0.79333), f32(-0.180868),
				f32(0.128495)],
			[f32(0.816108), f32(0.691169), f32(-0.130218)],
			[f32(0.85513), f32(-0.494777),
				f32(-0.42971)],
			[f32(0.992854), f32(0.132827), f32(-0.396611)]]
		faces:    [[9, 11, 18], [16, 23, 25], [10, 19, 12], [3, 6, 1],
			[2, 0, 4], [17, 13, 7], [15, 5, 8], [21, 14, 22],
			[26, 28, 29], [24, 27, 20], [19, 22, 12], [12, 22, 14],
			[12, 14, 6], [6, 14, 8], [6, 8, 1], [1, 8, 5], [1, 5, 0],
			[0, 5, 7], [0, 7, 4], [4, 7, 13], [4, 13, 11], [11, 13, 20],
			[11, 20, 18], [18, 20, 27], [18, 27, 23], [23, 27, 29],
			[23, 29, 25], [25, 29, 28], [25, 28, 19], [19, 28, 22],
			[9, 2, 4, 11], [16, 9, 18, 23], [10, 16, 25, 19],
			[3, 10, 12, 6], [2, 3, 1, 0], [17, 24, 20, 13], [15, 17, 7, 5],
			[21, 15, 8, 14], [26, 21, 22, 28], [24, 26, 29, 27],
			[2, 9, 16, 10, 3], [24, 17, 15, 21, 26]]
	},
	&Polyhedron{
		name:     'j47'
		vertexes: [[f32(-0.908535), f32(-0.523787), f32(-0.144699)],
			[f32(-0.894854), f32(-0.367641), f32(0.429886)],
			[f32(-0.853258), f32(0.048135),
				f32(-0.301436)],
			[f32(-0.839577), f32(0.20428), f32(0.273149)],
			[f32(-0.708763), f32(-0.381742),
				f32(-0.687498)],
			[f32(-0.672946), f32(0.027052), f32(0.816785)],
			[f32(-0.520247), f32(-0.782937),
				f32(0.225153)],
			[f32(-0.51634), f32(0.434114), f32(-0.605119)],
			[f32(-0.494204), f32(0.686763),
				f32(0.324579)],
			[f32(-0.422413), f32(-0.79035), f32(-0.362291)],
			[f32(-0.396391), f32(-0.493344),
				f32(0.730635)],
			[f32(-0.371845), f32(0.004237), f32(-0.991181)],
			[f32(-0.327573), f32(0.509534),
				f32(0.868216)],
			[f32(-0.294432), f32(0.828807), f32(-0.218221)],
			[f32(-0.140258), f32(-0.512752),
				f32(-0.807313)],
			[f32(-0.098153), f32(-0.032185), f32(0.961078)],
			[f32(-0.026471), f32(0.486719),
				f32(-0.939751)],
			[f32(-0.010949), f32(-1.00522), f32(0.010862)],
			[f32(0.009345), f32(0.895513),
				f32(0.564533)],
			[f32(0.189455), f32(-0.536653), f32(0.828749)],
			[f32(0.195436), f32(0.881412),
				f32(-0.552852)],
			[f32(0.209117), f32(1.03756), f32(0.021734)],
			[f32(0.218444), f32(-0.056175),
				f32(-0.93993)],
			[f32(0.260549), f32(0.424392), f32(0.828462)],
			[f32(0.427671), f32(-0.853012),
				f32(0.383905)],
			[f32(0.445587), f32(-0.556061), f32(-0.709199)],
			[f32(0.516681), f32(0.404984),
				f32(-0.709486)],
			[f32(0.525505), f32(-0.860425), f32(-0.203539)],
			[f32(0.542703), f32(0.70199),
				f32(0.38344)],
			[f32(0.640537), f32(0.694577),
				f32(-0.204005)],
			[f32(0.725908), f32(-0.391854), f32(0.614349)],
			[f32(0.769847), f32(0.202104),
				f32(0.614171)],
			[f32(0.884207), f32(-0.403849), f32(-0.336156)],
			[f32(0.928145), f32(0.190109),
				f32(-0.336334)],
			[f32(1.00806), f32(-0.114255), f32(0.169326)]]
		faces:    [[8, 12, 18], [13, 21, 20], [7, 16, 11], [2, 4, 0],
			[3, 1, 5], [30, 19, 24], [19, 15, 10], [24, 17, 27],
			[17, 6, 9], [27, 25, 32], [25, 14, 22], [32, 33, 34],
			[33, 26, 29], [34, 31, 30], [31, 28, 23], [16, 22, 11],
			[11, 22, 14], [11, 14, 4], [4, 14, 9], [4, 9, 0],
			[0, 9, 6], [0, 6, 1], [1, 6, 10], [1, 10, 5], [5, 10, 15],
			[5, 15, 12], [12, 15, 23], [12, 23, 18], [18, 23, 28],
			[18, 28, 21], [21, 28, 29], [21, 29, 20], [20, 29, 26],
			[20, 26, 16], [16, 26, 22], [8, 3, 5, 12], [13, 8, 18, 21],
			[7, 13, 20, 16], [2, 7, 11, 4], [3, 2, 0, 1], [3, 8, 13, 7, 2],
			[30, 24, 27, 32, 34], [30, 31, 23, 15, 19], [24, 19, 10, 6, 17],
			[27, 17, 9, 14, 25], [32, 25, 22, 26, 33], [34, 33, 29, 28, 31]]
	},
	&Polyhedron{
		name:     'j48'
		vertexes: [[f32(-1.02384), f32(0.34935), f32(0.211966)],
			[f32(-1.02284), f32(0.245289), f32(-0.329944)],
			[f32(-0.984402), f32(-0.132386),
				f32(0.478181)],
			[f32(-0.982778), f32(-0.300762), f32(-0.398647)],
			[f32(-0.959023), f32(-0.534178), f32(0.100801)],
			[f32(-0.762835), f32(0.690856),
				f32(-0.134076)],
			[f32(-0.724398), f32(0.313181), f32(0.674049)],
			[f32(-0.72177), f32(0.040743),
				f32(-0.74469)],
			[f32(-0.659577), f32(-0.570348), f32(0.562884)],
			[f32(-0.657953), f32(-0.738723),
				f32(-0.313945)],
			[f32(-0.302078), f32(0.865747), f32(0.11414)],
			[f32(-0.301074), f32(0.761686),
				f32(-0.427769)],
			[f32(-0.278322), f32(0.632332), f32(0.613589)],
			[f32(-0.275694), f32(0.359894),
				f32(-0.805149)],
			[f32(-0.238881), f32(0.150594), f32(0.879804)],
			[f32(-0.235633), f32(-0.186157),
				f32(-0.873853)],
			[f32(-0.198819), f32(-0.395456), f32(0.8111)],
			[f32(-0.196192), f32(-0.667893),
				f32(-0.607638)],
			[f32(-0.173439), f32(-0.797247), f32(0.43372)],
			[f32(-0.172436), f32(-0.901309),
				f32(-0.10819)],
			[f32(0.169627), f32(0.892069), f32(-0.170988)],
			[f32(0.181588), f32(0.824063),
				f32(0.376487)],
			[f32(0.183498), f32(0.626126), f32(-0.654287)],
			[f32(0.214813), f32(0.448086),
				f32(0.77902)],
			[f32(0.217902), f32(0.127816), f32(-0.888807)],
			[f32(0.25661), f32(-0.092255),
				f32(0.882858)],
			[f32(0.259699), f32(-0.412524), f32(-0.784969)],
			[f32(0.291015), f32(-0.590564),
				f32(0.648338)],
			[f32(0.292924), f32(-0.788502), f32(-0.382436)],
			[f32(0.304885), f32(-0.856507),
				f32(0.165038)],
			[f32(0.65102), f32(0.715912), f32(-0.375257)],
			[f32(0.670374), f32(0.605876),
				f32(0.510575)],
			[f32(0.706688), f32(-0.090371), f32(-0.754719)],
			[f32(0.738003), f32(-0.268411),
				f32(0.678589)],
			[f32(0.760446), f32(-0.698716), f32(-0.103406)],
			[f32(0.960498), f32(0.539035),
				f32(0.045972)],
			[f32(0.974369), f32(0.273093), f32(-0.437327)],
			[f32(0.993723), f32(0.163058),
				f32(0.448505)],
			[f32(1.01617), f32(-0.267247), f32(-0.333489)],
			[f32(1.02813), f32(-0.335253),
				f32(0.213985)]]
		faces:    [[0, 5, 1], [5, 10, 11], [1, 7, 3], [7, 13, 15],
			[3, 9, 4], [9, 17, 19], [4, 8, 2], [8, 18, 16], [2, 6, 0],
			[6, 14, 12], [35, 31, 37], [31, 21, 23], [37, 33, 39],
			[33, 25, 27], [39, 34, 38], [34, 29, 28], [38, 32, 36],
			[32, 26, 24], [36, 30, 35], [30, 22, 20], [17, 28, 19],
			[19, 28, 29], [19, 29, 18], [18, 29, 27], [18, 27, 16],
			[16, 27, 25], [16, 25, 14], [14, 25, 23], [14, 23, 12],
			[12, 23, 21], [12, 21, 10], [10, 21, 20], [10, 20, 11],
			[11, 20, 22], [11, 22, 13], [13, 22, 24], [13, 24, 15],
			[15, 24, 26], [15, 26, 17], [17, 26, 28], [0, 1, 3, 4, 2],
			[0, 6, 12, 10, 5], [1, 5, 11, 13, 7], [3, 7, 15, 17, 9],
			[4, 9, 19, 18, 8], [2, 8, 16, 14, 6], [35, 37, 39, 38, 36],
			[35, 30, 20, 21, 31], [37, 31, 23, 25, 33], [39, 33, 27, 29, 34],
			[38, 34, 28, 26, 32], [36, 32, 24, 22, 30]]
	},
	&Polyhedron{
		name:     'j49'
		vertexes: [[f32(-0.87547), f32(-0.255205), f32(-0.086794)],
			[f32(-0.276612), f32(-0.313401), f32(1.02999)],
			[f32(-0.236035), f32(0.801921),
				f32(-0.374595)],
			[f32(-0.051128), f32(-0.255205), f32(-1.05099)],
			[f32(0.218493), f32(-0.889481),
				f32(0.014004)],
			[f32(0.362823), f32(0.743725), f32(0.742188)],
			[f32(0.857929), f32(0.167645),
				f32(-0.273797)]]
		faces:    [[6, 3, 2], [3, 0, 2], [0, 3, 4], [2, 5, 6],
			[1, 0, 4], [6, 4, 3], [2, 0, 1, 5], [5, 1, 4, 6]]
	},
	&Polyhedron{
		name:     'j50'
		vertexes: [[f32(-0.878027), f32(-0.44614), f32(0.176652)],
			[f32(-0.85656), f32(0.548188), f32(-0.533)],
			[f32(-0.47761), f32(0.616903), f32(0.626496)],
			[f32(-0.069889), f32(-0.364329),
				f32(-0.736024)],
			[f32(0.239836), f32(-0.921955), f32(0.306031)],
			[f32(0.330528), f32(0.698715),
				f32(-0.286179)],
			[f32(0.640253), f32(0.141088), f32(0.755876)],
			[f32(1.07147), f32(-0.272471),
				f32(-0.309853)]]
		faces:    [[3, 0, 1], [1, 0, 2], [1, 2, 5], [4, 0, 3],
			[2, 6, 5], [4, 3, 7], [4, 7, 6], [6, 7, 5], [7, 3, 5],
			[1, 5, 3], [0, 4, 6, 2]]
	},
	&Polyhedron{
		name:     'j51'
		vertexes: [[f32(-0.837735), f32(-0.140456), f32(-0.298855)],
			[f32(-0.67808), f32(0.951266), f32(0.116678)],
			[f32(-0.424767), f32(0.019903),
				f32(0.793738)],
			[f32(-0.041529), f32(-0.887587), f32(0.145967)],
			[f32(-0.017092), f32(-0.613922),
				f32(-1.00056)],
			[f32(0.031619), f32(0.531638), f32(-0.726088)],
			[f32(0.444587), f32(0.691997),
				f32(0.366504)],
			[f32(0.695172), f32(-0.337344), f32(0.883883)],
			[f32(0.827825), f32(-0.215493),
				f32(-0.281266)]]
		faces:    [[1, 5, 0], [8, 4, 5], [4, 0, 5], [4, 3, 0],
			[8, 3, 4], [5, 6, 8], [8, 6, 7], [8, 7, 3], [3, 7, 2],
			[7, 6, 2], [3, 2, 0], [0, 2, 1], [2, 6, 1], [1, 6, 5]]
	},
	&Polyhedron{
		name:     'j52'
		vertexes: [[f32(-0.81481), f32(0.221521), f32(-0.662951)],
			[f32(-0.660297), f32(-0.683519), f32(-0.326712)],
			[f32(-0.53073), f32(0.852939), f32(0.027439)],
			[f32(-0.280723), f32(-0.611446),
				f32(0.571485)],
			[f32(-0.200646), f32(0.338137), f32(0.790362)],
			[f32(0.085423), f32(0.233517),
				f32(-1.04435)],
			[f32(0.239936), f32(-0.671523), f32(-0.708109)],
			[f32(0.369503), f32(0.864935),
				f32(-0.353959)],
			[f32(0.473247), f32(-0.295241), f32(1.10774)],
			[f32(0.619511), f32(-0.59945),
				f32(0.190087)],
			[f32(0.699587), f32(0.350133), f32(0.408964)]]
		faces:    [[3, 8, 4], [3, 9, 8], [4, 8, 10], [10, 8, 9],
			[1, 0, 5, 6], [3, 1, 6, 9], [2, 4, 10, 7], [0, 2, 7, 5],
			[0, 1, 3, 4, 2], [7, 10, 9, 6, 5]]
	},
	&Polyhedron{
		name:     'j53'
		vertexes: [[f32(-0.736376), f32(0.261231), f32(-0.409511)],
			[f32(-0.572247), f32(-0.640818), f32(-0.200191)],
			[f32(-0.430826), f32(0.786388), f32(0.30833)],
			[f32(-0.352398), f32(1.10393),
				f32(-0.573408)],
			[f32(-0.16526), f32(-0.673158), f32(0.647018)],
			[f32(-0.077857), f32(0.208904),
				f32(0.961301)],
			[f32(0.083202), f32(-1.29012), f32(-0.017868)],
			[f32(0.11049), f32(0.32145),
				f32(-0.814035)],
			[f32(0.274618), f32(-0.5806), f32(-0.604714)],
			[f32(0.416039), f32(0.846607),
				f32(-0.096194)],
			[f32(0.681606), f32(-0.61294), f32(0.242494)],
			[f32(0.769009), f32(0.269122),
				f32(0.556777)]]
		faces:    [[2, 3, 0], [2, 9, 3], [0, 3, 7], [7, 3, 9],
			[1, 6, 4], [1, 8, 6], [4, 6, 10], [10, 6, 8], [5, 4, 10, 11],
			[2, 5, 11, 9], [1, 0, 7, 8], [4, 5, 2, 0, 1], [8, 7, 9, 11, 10]]
	},
	&Polyhedron{
		name:     'j54'
		vertexes: [[f32(-0.973522), f32(0.38842), f32(-0.100967)],
			[f32(-0.837708), f32(-0.464036), f32(-0.18462)],
			[f32(-0.457167), f32(0.537479),
				f32(-0.781617)],
			[f32(-0.449574), f32(0.863826), f32(0.400622)],
			[f32(-0.321353), f32(-0.314977),
				f32(-0.865269)],
			[f32(-0.177946), f32(-0.841086), f32(0.233318)],
			[f32(0.066781), f32(1.01288),
				f32(-0.280028)],
			[f32(0.210188), f32(0.486776), f32(0.818559)],
			[f32(0.338409), f32(-0.692027),
				f32(-0.447332)],
			[f32(0.346002), f32(-0.365679), f32(0.734907)],
			[f32(0.666998), f32(-1.0308),
				f32(0.280259)],
			[f32(0.726543), f32(0.635835), f32(0.13791)],
			[f32(0.862357), f32(-0.216621),
				f32(0.054258)]]
		faces:    [[5, 10, 9], [5, 8, 10], [9, 10, 12], [12, 10, 8],
			[1, 0, 2, 4], [5, 1, 4, 8], [7, 9, 12, 11], [3, 7, 11, 6],
			[0, 3, 6, 2], [0, 1, 5, 9, 7, 3], [11, 12, 8, 4, 2, 6]]
	},
	&Polyhedron{
		name:     'j55'
		vertexes: [[f32(-1.12956), f32(0.266324), f32(0.624401)],
			[f32(-0.925111), f32(0.008507), f32(-0.145991)],
			[f32(-0.655368), f32(-0.416841),
				f32(0.523404)],
			[f32(-0.5883), f32(0.71007), f32(0.164074)],
			[f32(-0.438148), f32(0.074567),
				f32(-0.824427)],
			[f32(-0.318557), f32(0.284721), f32(0.83347)],
			[f32(-0.101337), f32(0.77613),
				f32(-0.514362)],
			[f32(0.101337), f32(-0.77613), f32(0.514363)],
			[f32(0.318557), f32(-0.284721),
				f32(-0.833468)],
			[f32(0.438148), f32(-0.074567), f32(0.824429)],
			[f32(0.5883), f32(-0.710069),
				f32(-0.164073)],
			[f32(0.655368), f32(0.416842), f32(-0.523403)],
			[f32(0.925111), f32(-0.008507),
				f32(0.145993)],
			[f32(1.12956), f32(-0.266324), f32(-0.624399)]]
		faces:    [[12, 13, 11], [12, 10, 13], [11, 13, 8], [8, 13, 10],
			[3, 0, 5], [3, 1, 0], [5, 0, 2], [2, 0, 1], [9, 5, 2, 7],
			[12, 9, 7, 10], [6, 11, 8, 4], [3, 6, 4, 1], [5, 9, 12, 11, 6, 3],
			[4, 8, 10, 7, 2, 1]]
	},
	&Polyhedron{
		name:     'j56'
		vertexes: [[f32(-1.11176), f32(0.435562), f32(-0.458586)],
			[f32(-0.808867), f32(0.159752), f32(0.27642)],
			[f32(-0.700013), f32(-0.297342),
				f32(-0.421621)],
			[f32(-0.454926), f32(0.822531), f32(-0.102389)],
			[f32(-0.346072), f32(0.365437),
				f32(-0.80043)],
			[f32(-0.331474), f32(-0.383478), f32(0.706586)],
			[f32(-0.22262), f32(-0.840572),
				f32(0.008545)],
			[f32(0.189019), f32(-1.0446), f32(0.713507)],
			[f32(0.376408), f32(0.942079),
				f32(-0.051032)],
			[f32(0.485263), f32(0.484985), f32(-0.749073)],
			[f32(0.49986), f32(-0.26393),
				f32(0.757943)],
			[f32(0.608714), f32(-0.721024), f32(0.059902)],
			[f32(0.853802), f32(0.398849),
				f32(0.379134)],
			[f32(0.962656), f32(-0.058246), f32(-0.318907)]]
		faces:    [[3, 0, 1], [3, 4, 0], [1, 0, 2], [2, 0, 4],
			[5, 7, 10], [5, 6, 7], [10, 7, 11], [11, 7, 6], [8, 12, 13, 9],
			[3, 8, 9, 4], [5, 1, 2, 6], [12, 10, 11, 13], [12, 8, 3, 1, 5, 10],
			[6, 2, 4, 9, 13, 11]]
	},
	&Polyhedron{
		name:     'j57'
		vertexes: [[f32(-0.902174), f32(-0.044182), f32(-0.142406)],
			[f32(-0.852256), f32(-0.16038), f32(-0.950443)],
			[f32(-0.65694), f32(0.352221),
				f32(0.529639)],
			[f32(-0.484062), f32(0.483825), f32(-0.606421)],
			[f32(-0.454289), f32(-0.660407),
				f32(-0.440037)],
			[f32(-0.238829), f32(0.880229), f32(0.065624)],
			[f32(-0.184058), f32(0.919718),
				f32(0.880707)],
			[f32(-0.036177), f32(-0.1324), f32(-0.904053)],
			[f32(0.036178), f32(0.1324), f32(0.904052)],
			[f32(0.238829), f32(-0.880229),
				f32(-0.065625)],
			[f32(0.454289), f32(0.660407), f32(0.440037)],
			[f32(0.484063), f32(-0.483825),
				f32(0.60642)],
			[f32(0.656941), f32(-0.352221), f32(-0.52964)],
			[f32(0.902174), f32(0.044182),
				f32(0.142405)],
			[f32(1.03631), f32(-0.759338), f32(0.069736)]]
		faces:    [[9, 14, 11], [9, 12, 14], [11, 14, 13], [13, 14, 12],
			[8, 6, 2], [8, 10, 6], [2, 6, 5], [5, 6, 10], [0, 1, 4],
			[0, 3, 1], [4, 1, 7], [7, 1, 3], [9, 4, 7, 12], [8, 11, 13, 10],
			[0, 2, 5, 3], [0, 4, 9, 11, 8, 2], [10, 13, 12, 7, 3, 5]]
	},
	&Polyhedron{
		name:     'j58'
		vertexes: [[f32(-0.906673), f32(0.136106), f32(0.246909)],
			[f32(-0.827056), f32(0.097501), f32(-0.456089)],
			[f32(-0.822039), f32(0.728118),
				f32(-0.133084)],
			[f32(-0.682157), f32(-0.474972), f32(0.526574)],
			[f32(-0.553334), f32(-0.537436),
				f32(-0.610901)],
			[f32(-0.48677), f32(0.654002), f32(0.486704)],
			[f32(-0.463781), f32(-0.891244),
				f32(-0.003583)],
			[f32(-0.357947), f32(0.591537), f32(-0.650771)],
			[f32(-0.147639), f32(0.935474),
				f32(-0.068093)],
			[f32(-0.123496), f32(-0.334743), f32(0.939211)],
			[f32(-0.00274), f32(0.363001),
				f32(0.91457)],
			[f32(0.084945), f32(-0.435813), f32(-0.901263)],
			[f32(0.2057), f32(0.261931),
				f32(-0.925903)],
			[f32(0.229843), f32(-1.00829), f32(0.0814)],
			[f32(0.440151), f32(-0.664349), f32(0.664079)],
			[f32(0.545986), f32(0.818432),
				f32(0.01689)],
			[f32(0.568974), f32(-0.726814), f32(-0.473396)],
			[f32(0.635538), f32(0.464625),
				f32(0.624209)],
			[f32(0.764361), f32(0.40216), f32(-0.513266)],
			[f32(0.90926), f32(-0.170313),
				f32(0.469397)],
			[f32(0.988877), f32(-0.208918), f32(-0.233601)]]
		faces:    [[2, 0, 5], [2, 5, 8], [2, 1, 0], [2, 7, 1],
			[7, 2, 8], [18, 20, 16, 11, 12], [6, 4, 11, 16, 13],
			[1, 7, 12, 11, 4], [8, 15, 18, 12, 7], [17, 19, 20, 18, 15],
			[14, 13, 16, 20, 19], [19, 17, 10, 9, 14], [15, 8, 5, 10, 17],
			[4, 6, 3, 0, 1], [13, 14, 9, 3, 6], [3, 9, 10, 5, 0]]
	},
	&Polyhedron{
		name:     'j59'
		vertexes: [[f32(-0.987924), f32(-0.168105), f32(-0.565605)],
			[f32(-0.950092), f32(-0.216897), f32(0.133657)],
			[f32(-0.877263), f32(0.407337),
				f32(-0.179083)],
			[f32(-0.637339), f32(-0.699196), f32(-0.269274)],
			[f32(-0.609869), f32(-0.193139), f32(0.747222)],
			[f32(-0.519498), f32(0.310837),
				f32(-0.775297)],
			[f32(-0.492028), f32(0.816894), f32(0.241199)],
			[f32(-0.371218), f32(-0.373038),
				f32(-0.831038)],
			[f32(-0.32677), f32(0.445779), f32(0.813687)],
			[f32(-0.103824), f32(-0.973514),
				f32(0.095267)],
			[f32(-0.086847), f32(-0.660753), f32(0.723496)],
			[f32(0.086847), f32(0.660753),
				f32(-0.723496)],
			[f32(0.103824), f32(0.973513), f32(-0.095267)],
			[f32(0.32677), f32(-0.44578),
				f32(-0.813687)],
			[f32(0.371218), f32(0.373038), f32(0.831038)],
			[f32(0.492028), f32(-0.816894),
				f32(-0.241199)],
			[f32(0.519498), f32(-0.310837), f32(0.775297)],
			[f32(0.609869), f32(0.193139),
				f32(-0.747222)],
			[f32(0.637339), f32(0.699195), f32(0.269274)],
			[f32(0.877262), f32(-0.407338),
				f32(0.179083)],
			[f32(0.950092), f32(0.216897), f32(-0.133657)],
			[f32(0.987924), f32(0.168105),
				f32(0.565605)]]
		faces:    [[0, 7, 3], [0, 3, 1], [0, 5, 7], [0, 2, 5],
			[2, 0, 1], [21, 18, 14], [21, 14, 16], [21, 20, 18],
			[21, 19, 20], [19, 21, 16], [6, 8, 14, 18, 12], [17, 11, 12, 18, 20],
			[5, 2, 6, 12, 11], [1, 4, 8, 6, 2], [10, 16, 14, 8, 4],
			[4, 1, 3, 9, 10], [11, 17, 13, 7, 5], [20, 19, 15, 13, 17],
			[16, 10, 9, 15, 19], [15, 9, 3, 7, 13]]
	},
	&Polyhedron{
		name:     'j60'
		vertexes: [[f32(-0.858966), f32(-0.256781), f32(-0.362035)],
			[f32(-0.807204), f32(-0.391109), f32(0.326114)],
			[f32(-0.719263), f32(0.425042),
				f32(-0.461407)],
			[f32(-0.63551), f32(0.207695), f32(0.652043)],
			[f32(-0.58116), f32(0.712103),
				f32(0.165328)],
			[f32(-0.46306), f32(-0.410585), f32(0.938862)],
			[f32(-0.364654), f32(-0.630479),
				f32(-0.694119)],
			[f32(-0.311484), f32(0.996138), f32(-0.418515)],
			[f32(-0.280902), f32(-0.847826),
				f32(0.419331)],
			[f32(-0.13861), f32(0.472734), f32(-0.854906)],
			[f32(-0.007391), f32(-0.995764),
				f32(-0.211209)],
			[f32(-0.003096), f32(0.121058), f32(0.946694)],
			[f32(0.08055), f32(-0.179614),
				f32(-0.99873)],
			[f32(0.084846), f32(0.937209), f32(0.159173)],
			[f32(0.216065), f32(-0.531289),
				f32(0.80287)],
			[f32(0.358357), f32(0.789271), f32(-0.471366)],
			[f32(0.442109), f32(0.571923),
				f32(0.642084)],
			[f32(0.658614), f32(-0.770659), f32(-0.217364)],
			[f32(0.712965), f32(-0.26625),
				f32(-0.704079)],
			[f32(0.796718), f32(-0.483597), f32(0.409371)],
			[f32(0.884659), f32(0.332554),
				f32(-0.37815)],
			[f32(0.936421), f32(0.198226), f32(0.31)]]
		faces:    [[7, 13, 15], [7, 15, 9], [7, 4, 13], [7, 2, 4],
			[2, 7, 9], [5, 1, 8], [5, 8, 14], [5, 3, 1], [5, 11, 3],
			[11, 5, 14], [0, 6, 10, 8, 1], [19, 14, 8, 10, 17],
			[4, 2, 0, 1, 3], [9, 12, 6, 0, 2], [18, 17, 10, 6, 12],
			[12, 9, 15, 20, 18], [3, 11, 16, 13, 4], [14, 19, 21, 16, 11],
			[17, 18, 20, 21, 19], [21, 20, 15, 13, 16]]
	},
	&Polyhedron{
		name:     'j61'
		vertexes: [[f32(-0.875027), f32(-0.215344), f32(-0.354115)],
			[f32(-0.822602), f32(-0.401147), f32(0.315989)],
			[f32(-0.733096), f32(0.465836),
				f32(-0.400606)],
			[f32(-0.648272), f32(0.1652), f32(0.683645)],
			[f32(-0.625957), f32(0.049095),
				f32(-0.949385)],
			[f32(-0.592955), f32(0.701024), f32(0.240765)],
			[f32(-0.479753), f32(-0.469083),
				f32(0.919437)],
			[f32(-0.387571), f32(-0.561993), f32(-0.712628)],
			[f32(-0.302747), f32(-0.862629), f32(0.371622)],
			[f32(-0.157924), f32(0.540178),
				f32(-0.787852)],
			[f32(-0.033883), f32(-0.962037), f32(-0.264098)],
			[f32(-0.020675), f32(0.053739), f32(0.966503)],
			[f32(0.055623), f32(-0.095055),
				f32(-0.980693)],
			[f32(0.068831), f32(0.920721), f32(0.249908)],
			[f32(0.192872), f32(-0.581494),
				f32(0.773662)],
			[f32(0.337694), f32(0.821313), f32(-0.385812)],
			[f32(0.422519), f32(0.520677),
				f32(0.698439)],
			[f32(0.627903), f32(-0.74234), f32(-0.254955)],
			[f32(0.683221), f32(-0.206515),
				f32(-0.697835)],
			[f32(0.756251), f32(0.83314), f32(0.171845)],
			[f32(0.768045), f32(-0.507151),
				f32(0.386416)],
			[f32(0.85755), f32(0.359831), f32(-0.330178)],
			[f32(0.909975), f32(0.174028),
				f32(0.339925)]]
		faces:    [[6, 3, 1], [6, 1, 8], [6, 11, 3], [6, 14, 11],
			[14, 6, 8], [19, 22, 21], [19, 21, 15], [19, 16, 22],
			[19, 13, 16], [13, 19, 15], [4, 0, 2], [4, 2, 9],
			[4, 7, 0], [4, 12, 7], [12, 4, 9], [20, 17, 18, 21, 22],
			[9, 15, 21, 18, 12], [11, 14, 20, 22, 16], [8, 10, 17, 20, 14],
			[7, 12, 18, 17, 10], [10, 8, 1, 0, 7], [16, 13, 5, 3, 11],
			[15, 9, 2, 5, 13], [2, 0, 1, 3, 5]]
	},
	&Polyhedron{
		name:     'j62'
		vertexes: [[f32(-0.821855), f32(0.223834), f32(-0.340481)],
			[f32(-0.71039), f32(-0.701977), f32(0.157898)],
			[f32(-0.692806), f32(0.20039),
				f32(0.708676)],
			[f32(-0.215696), f32(-0.533443), f32(-0.761235)],
			[f32(-0.187244), f32(0.926618), f32(0.129942)],
			[f32(-0.006891), f32(-0.571377),
				f32(0.936336)],
			[f32(0.107626), f32(0.473083), f32(-0.778513)],
			[f32(0.793541), f32(-0.298683),
				f32(-0.550854)],
			[f32(0.811125), f32(0.603684), f32(-7.6e-05)],
			[f32(0.92259), f32(-0.322128),
				f32(0.498303)]]
		faces:    [[6, 3, 0], [0, 3, 1], [1, 5, 2], [1, 2, 0],
			[2, 4, 0], [4, 8, 6], [4, 6, 0], [9, 7, 8], [7, 6, 8],
			[7, 3, 6], [1, 3, 7, 9, 5], [2, 5, 9, 8, 4]]
	},
	&Polyhedron{
		name:     'j63'
		vertexes: [[f32(-0.799898), f32(0.494585), f32(-0.153719)],
			[f32(-0.680241), f32(-0.086273), f32(0.717027)],
			[f32(-0.306176), f32(0.002547),
				f32(-0.943688)],
			[f32(-0.112567), f32(-0.9373), f32(0.465209)],
			[f32(-0.077419), f32(0.764103),
				f32(0.564122)],
			[f32(0.118618), f32(-0.882406), f32(-0.56117)],
			[f32(0.153766), f32(0.818996),
				f32(-0.462256)],
			[f32(0.841097), f32(-0.612888), f32(0.156672)],
			[f32(0.86282), f32(0.438637),
				f32(0.217804)]]
		faces:    [[0, 4, 6], [4, 8, 6], [6, 2, 0], [0, 1, 4],
			[5, 7, 3], [6, 8, 7, 5, 2], [0, 2, 5, 3, 1], [7, 8, 4, 1, 3]]
	},
	&Polyhedron{
		name:     'j64'
		vertexes: [[f32(-0.777985), f32(-0.188235), f32(-0.285228)],
			[f32(-0.489362), f32(-0.260552), f32(0.643961)],
			[f32(-0.32442), f32(0.578558),
				f32(-0.683014)],
			[f32(-0.099589), f32(-0.843165), f32(-0.034687)],
			[f32(0.142581), f32(0.461547), f32(0.820446)],
			[f32(0.24452), f32(0.980145), f32(0.00033)],
			[f32(0.634293), f32(0.397531), f32(-0.678318)],
			[f32(0.773247), f32(-0.481142),
				f32(-0.27763)],
			[f32(0.922916), f32(0.325215), f32(0.250871)],
			[f32(-1.0262), f32(-0.969903), f32(0.24327)]]
		faces:    [[6, 5, 8], [5, 4, 8], [8, 7, 6], [6, 2, 5],
			[9, 1, 0], [9, 0, 3], [9, 3, 1], [8, 4, 1, 3, 7],
			[6, 7, 3, 0, 2], [1, 4, 5, 2, 0]]
	},
	&Polyhedron{
		name:     'j65'
		vertexes: [[f32(-0.91403), f32(0.409064), f32(-0.602734)],
			[f32(-0.830829), f32(0.815648), f32(0.102539)],
			[f32(-0.699591), f32(-0.379344),
				f32(-0.648261)],
			[f32(-0.533188), f32(0.433825), f32(0.762285)],
			[f32(-0.401951), f32(-0.761167),
				f32(0.011485)],
			[f32(-0.338469), f32(0.986004), f32(-0.528495)],
			[f32(-0.318749), f32(-0.354582),
				f32(0.716757)],
			[f32(0.090409), f32(-0.59081), f32(-0.619549)],
			[f32(0.251663), f32(-0.893891),
				f32(0.485632)],
			[f32(0.256812), f32(0.222359), f32(0.790997)],
			[f32(0.451531), f32(0.774538),
				f32(-0.499782)],
			[f32(0.66597), f32(-0.013869), f32(-0.545309)],
			[f32(0.744023), f32(-0.723534),
				f32(-0.145401)],
			[f32(0.749172), f32(0.392715), f32(0.159963)],
			[f32(0.827225), f32(-0.31695),
				f32(0.559871)]]
		faces:    [[12, 7, 11], [10, 13, 11], [14, 13, 9], [9, 3, 6],
			[0, 1, 5], [4, 2, 7], [6, 4, 8], [14, 8, 12], [12, 8, 4, 7],
			[13, 14, 12, 11], [14, 9, 6, 8], [11, 7, 2, 0, 5, 10],
			[13, 10, 5, 1, 3, 9], [3, 1, 0, 2, 4, 6]]
	},
	&Polyhedron{
		name:     'j66'
		vertexes: [[f32(-0.935384), f32(0.507278), f32(-0.272116)],
			[f32(-0.915801), f32(0.536228), f32(0.283002)],
			[f32(-0.882043), f32(0.099694),
				f32(-0.646826)],
			[f32(-0.834764), f32(0.169584), f32(0.693348)],
			[f32(-0.787023), f32(-0.447768),
				f32(-0.621628)],
			[f32(-0.739744), f32(-0.377878), f32(0.718546)],
			[f32(-0.705986), f32(-0.814411),
				f32(-0.211282)],
			[f32(-0.686402), f32(-0.785462), f32(0.343836)],
			[f32(-0.561956), f32(0.553237),
				f32(-0.681771)],
			[f32(-0.514677), f32(0.623127), f32(0.658404)],
			[f32(-0.332557), f32(-0.768453),
				f32(-0.620937)],
			[f32(-0.285278), f32(-0.698562), f32(0.719237)],
			[f32(-0.014265), f32(0.647182),
				f32(-0.705992)],
			[f32(0.033015), f32(0.717073), f32(0.634183)],
			[f32(0.215134), f32(-0.674508),
				f32(-0.645158)],
			[f32(0.262413), f32(-0.604617), f32(0.695016)],
			[f32(0.386859), f32(0.734081),
				f32(-0.330591)],
			[f32(0.406443), f32(0.763031), f32(0.224528)],
			[f32(0.440201), f32(0.326497),
				f32(-0.705301)],
			[f32(0.48748), f32(0.396388), f32(0.634874)],
			[f32(0.535221), f32(-0.220964),
				f32(-0.680103)],
			[f32(0.5825), f32(-0.151074), f32(0.660072)],
			[f32(0.616258), f32(-0.587608),
				f32(-0.269757)],
			[f32(0.635842), f32(-0.558659), f32(0.285361)],
			[f32(0.831438), f32(0.541255),
				f32(-0.057559)],
			[f32(0.884779), f32(0.13367), f32(-0.432269)],
			[f32(0.912475), f32(0.174611),
				f32(0.352787)],
			[f32(0.965816), f32(-0.232973), f32(-0.021924)]]
		faces:    [[24, 16, 17], [26, 19, 21], [27, 23, 22], [25, 20, 18],
			[21, 15, 23], [5, 7, 11], [17, 13, 19], [1, 3, 9],
			[18, 12, 16], [2, 0, 8], [22, 14, 20], [6, 4, 10],
			[25, 24, 26, 27], [24, 25, 18, 16], [26, 24, 17, 19],
			[27, 26, 21, 23], [25, 27, 22, 20], [23, 15, 11, 7, 6, 10, 14, 22],
			[20, 14, 10, 4, 2, 8, 12, 18], [16, 12, 8, 0, 1, 9, 13, 17],
			[19, 13, 9, 3, 5, 11, 15, 21], [4, 6, 7, 5, 3, 1, 0, 2]]
	},
	&Polyhedron{
		name:     'j67'
		vertexes: [[f32(-0.85468), f32(-0.304544), f32(0.321795)],
			[f32(-0.813538), f32(0.214997), f32(0.467663)],
			[f32(-0.753988), f32(-0.584165),
				f32(-0.130495)],
			[f32(-0.662946), f32(-0.809677), f32(0.352981)],
			[f32(-0.654663), f32(0.670118),
				f32(0.221662)],
			[f32(-0.570447), f32(-0.460068), f32(-0.624262)],
			[f32(-0.567052), f32(-0.168344), f32(0.759532)],
			[f32(-0.471123), f32(0.794216),
				f32(-0.272106)],
			[f32(-0.411573), f32(-0.004947), f32(-0.870263)],
			[f32(-0.375319), f32(-0.673477), f32(0.790718)],
			[f32(-0.370431), f32(0.514594),
				f32(-0.724396)],
			[f32(-0.323962), f32(-0.84341), f32(-0.332393)],
			[f32(-0.23292), f32(-1.06892),
				f32(0.151083)],
			[f32(-0.183495), f32(0.930415), f32(0.165631)],
			[f32(-0.059594), f32(-0.25535),
				f32(0.926295)],
			[f32(-0.054707), f32(0.932721), f32(-0.588818)],
			[f32(0.054707), f32(-0.932721),
				f32(0.588819)],
			[f32(0.059595), f32(0.25535), f32(-0.926294)],
			[f32(0.183496), f32(-0.930415),
				f32(-0.16563)],
			[f32(0.23292), f32(1.06892), f32(-0.151082)],
			[f32(0.323962), f32(0.84341), f32(0.332394)],
			[f32(0.370432), f32(-0.514594),
				f32(0.724397)],
			[f32(0.37532), f32(0.673477), f32(-0.790717)],
			[f32(0.411574), f32(0.004947),
				f32(0.870264)],
			[f32(0.471123), f32(-0.794216), f32(0.272106)],
			[f32(0.567053), f32(0.168344),
				f32(-0.759531)],
			[f32(0.570448), f32(0.460068), f32(0.624263)],
			[f32(0.654664), f32(-0.670118),
				f32(-0.221661)],
			[f32(0.662947), f32(0.809677), f32(-0.35298)],
			[f32(0.753989), f32(0.584165),
				f32(0.130496)],
			[f32(0.813538), f32(-0.214997), f32(-0.467662)],
			[f32(0.85468), f32(0.304544),
				f32(-0.321795)]]
		faces:    [[22, 25, 17], [15, 10, 7], [19, 13, 20], [28, 29, 31],
			[9, 14, 6], [3, 0, 2], [12, 11, 18], [16, 24, 21],
			[7, 4, 13], [0, 6, 1], [17, 8, 10], [11, 2, 5], [31, 30, 25],
			[24, 18, 27], [20, 26, 29], [14, 21, 23], [28, 22, 15, 19],
			[22, 28, 31, 25], [15, 22, 17, 10], [19, 15, 7, 13],
			[28, 19, 20, 29], [16, 9, 3, 12], [9, 16, 21, 14],
			[3, 9, 6, 0], [12, 3, 2, 11], [16, 12, 18, 24], [13, 4, 1, 6, 14, 23, 26, 20],
			[29, 26, 23, 21, 24, 27, 30, 31], [25, 30, 27, 18, 11, 5, 8, 17],
			[10, 8, 5, 2, 0, 1, 4, 7]]
	},
	&Polyhedron{
		name:     'j68'
		vertexes: [[f32(-1.05373), f32(-0.062801), f32(0.140871)],
			[f32(-1.04773), f32(-0.006643), f32(-0.190675)],
			[f32(-0.967657), f32(0.064553),
				f32(0.440012)],
			[f32(-0.951944), f32(0.211579), f32(-0.427988)],
			[f32(-0.942283), f32(-0.266176),
				f32(0.38445)],
			[f32(-0.92657), f32(-0.11915), f32(-0.483549)],
			[f32(-0.822385), f32(0.326776),
				f32(0.592485)],
			[f32(-0.802963), f32(0.50851), f32(-0.480421)],
			[f32(-0.755954), f32(-0.539085),
				f32(0.447023)],
			[f32(-0.736532), f32(-0.35735), f32(-0.625883)],
			[f32(-0.673403), f32(0.623707),
				f32(0.540051)],
			[f32(-0.65769), f32(0.770733), f32(-0.327948)],
			[f32(-0.577618), f32(0.841928),
				f32(0.302738)],
			[f32(-0.571617), f32(0.898087), f32(-0.028808)],
			[f32(-0.565916), f32(-0.777285),
				f32(0.304689)],
			[f32(-0.561955), f32(0.420332), f32(0.78363)],
			[f32(-0.550203), f32(-0.630259),
				f32(-0.56331)],
			[f32(-0.536531), f32(0.658225), f32(-0.620822)],
			[f32(-0.479842), f32(-0.64993),
				f32(0.603829)],
			[f32(-0.454419), f32(-0.412037), f32(-0.800623)],
			[f32(-0.444757), f32(-0.889793), f32(0.011815)],
			[f32(-0.438755), f32(-0.833633),
				f32(-0.319731)],
			[f32(-0.311187), f32(0.991643), f32(0.162337)],
			[f32(-0.285843), f32(0.309485),
				f32(0.940436)],
			[f32(-0.254418), f32(0.603538), f32(-0.795562)],
			[f32(-0.219412), f32(-0.556374),
				f32(0.794974)],
			[f32(-0.187987), f32(-0.262321), f32(-0.941024)],
			[f32(-0.162643), f32(-0.944479), f32(-0.162925)],
			[f32(-0.099515), f32(0.036577), f32(1.00301)],
			[f32(-0.07414), f32(-0.294152),
				f32(0.947447)],
			[f32(-0.06438), f32(0.365339), f32(-0.937896)],
			[f32(-0.039006), f32(0.034609),
				f32(-0.993458)],
			[f32(0.024123), f32(1.01567), f32(0.172476)],
			[f32(0.049467), f32(0.333508), f32(0.950575)],
			[f32(0.080892), f32(0.627561),
				f32(-0.785423)],
			[f32(0.115898), f32(-0.532352), f32(0.805113)],
			[f32(0.147323), f32(-0.238299),
				f32(-0.930885)],
			[f32(0.172667), f32(-0.920457), f32(-0.152786)],
			[f32(0.300235), f32(0.90482),
				f32(0.329282)],
			[f32(0.306237), f32(0.960979), f32(-0.002264)],
			[f32(0.315898), f32(0.483223),
				f32(0.810173)],
			[f32(0.341322), f32(0.721117), f32(-0.594278)],
			[f32(0.398011), f32(-0.587039),
				f32(0.630373)],
			[f32(0.411683), f32(0.701445), f32(0.572861)],
			[f32(0.423435), f32(-0.349145),
				f32(-0.774079)],
			[f32(0.427396), f32(0.848471), f32(-0.295138)],
			[f32(0.433096), f32(-0.826901),
				f32(0.038358)],
			[f32(0.439098), f32(-0.770742), f32(-0.293188)],
			[f32(0.51917), f32(-0.699547),
				f32(0.337499)],
			[f32(0.534883), f32(-0.55252), f32(-0.5305)],
			[f32(0.598012), f32(0.428536), f32(0.635433)],
			[f32(0.617434), f32(0.610271),
				f32(-0.437472)],
			[f32(0.664443), f32(-0.437324), f32(0.489972)],
			[f32(0.683864), f32(-0.255589),
				f32(-0.582934)],
			[f32(0.721659), f32(-0.657508), f32(0.072275)],
			[f32(0.727661), f32(-0.601349),
				f32(-0.259271)],
			[f32(0.78805), f32(0.190336), f32(0.493099)],
			[f32(0.803762), f32(0.337363), f32(-0.3749)],
			[f32(0.813424), f32(-0.140393),
				f32(0.437538)],
			[f32(0.829136), f32(0.006634), f32(-0.430461)],
			[f32(0.866931), f32(-0.395285),
				f32(0.224748)],
			[f32(0.876642), f32(-0.304418), f32(-0.311705)],
			[f32(0.909209), f32(0.077829),
				f32(0.200225)],
			[f32(0.91521), f32(0.133987), f32(-0.131321)],
			[f32(0.962716), f32(-0.177064),
				f32(-0.012565)]]
		faces:    [[34, 30, 24], [45, 51, 41], [36, 26, 31], [53, 49, 44],
			[16, 9, 19], [27, 20, 21], [1, 3, 5], [4, 2, 0], [11, 17, 7],
			[12, 22, 13], [62, 56, 58], [59, 57, 63], [43, 40, 50],
			[39, 32, 38], [23, 28, 33], [10, 6, 15], [25, 35, 29],
			[8, 14, 18], [48, 52, 42], [47, 46, 37], [54, 48, 46],
			[55, 47, 49], [61, 53, 59], [62, 64, 63], [60, 58, 52],
			[54, 60, 52, 48], [55, 54, 46, 47], [61, 55, 49, 53],
			[64, 61, 59, 63], [60, 64, 62, 58], [60, 54, 55, 61, 64],
			[31, 26, 19, 9, 5, 3, 7, 17, 24, 30], [59, 53, 44, 36, 31, 30, 34, 41, 51, 57],
			[37, 27, 21, 16, 19, 26, 36, 44, 49, 47], [8, 4, 0, 1, 5, 9, 16, 21, 20, 14],
			[10, 12, 13, 11, 7, 3, 1, 0, 2, 6], [39, 45, 41, 34, 24, 17, 11, 13, 22, 32],
			[50, 40, 33, 28, 29, 35, 42, 52, 58, 56], [45, 39, 38, 43, 50, 56, 62, 63, 57, 51],
			[12, 10, 15, 23, 33, 40, 43, 38, 32, 22], [4, 8, 18, 25, 29, 28, 23, 15, 6, 2],
			[27, 37, 46, 48, 42, 35, 25, 18, 14, 20]]
	},
	&Polyhedron{
		name:     'j69'
		vertexes: [[f32(-0.988041), f32(0.082361), f32(-0.032394)],
			[f32(-0.940439), f32(0.10562), f32(0.297446)],
			[f32(-0.93903), f32(-0.112232),
				f32(-0.299475)],
			[f32(-0.911497), f32(0.377114), f32(0.10495)],
			[f32(-0.814408), f32(-0.051339),
				f32(0.564056)],
			[f32(-0.812127), f32(-0.403831), f32(-0.401783)],
			[f32(-0.783185), f32(-0.132338), f32(-0.594279)],
			[f32(-0.738637), f32(0.65944), f32(0.060095)],
			[f32(-0.658086), f32(-0.328563),
				f32(0.665601)],
			[f32(-0.655805), f32(-0.681055), f32(-0.300238)],
			[f32(-0.621075), f32(-0.575598), f32(-0.615315)],
			[f32(-0.592133), f32(-0.304105), f32(-0.807812)],
			[f32(-0.581542), f32(-0.03381), f32(0.802944)],
			[f32(-0.580033), f32(0.029724),
				f32(-0.8042)],
			[f32(-0.535485), f32(0.821501), f32(-0.149826)],
			[f32(-0.531183), f32(-0.620162),
				f32(0.563294)],
			[f32(-0.529773), f32(-0.838014), f32(-0.033627)],
			[f32(-0.487884), f32(0.844761), f32(0.180013)],
			[f32(-0.482172), f32(-0.814755),
				f32(0.296212)],
			[f32(-0.407173), f32(0.31205), f32(-0.849055)],
			[f32(-0.37964), f32(0.801396),
				f32(-0.44463)],
			[f32(-0.373928), f32(-0.858119), f32(-0.328432)],
			[f32(-0.339198), f32(-0.752663), f32(-0.643508)],
			[f32(-0.33079), f32(0.15151), f32(0.922864)],
			[f32(-0.330629), f32(0.606803),
				f32(-0.711711)],
			[f32(-0.292369), f32(-0.313377), f32(-0.954974)],
			[f32(-0.28027), f32(0.020452), f32(-0.951362)],
			[f32(-0.255019), f32(0.862289),
				f32(0.418901)],
			[f32(-0.249306), f32(-0.797226), f32(0.5351)],
			[f32(-0.157929), f32(0.433837),
				f32(0.878008)],
			[f32(-0.136047), f32(-0.590601), f32(-0.85343)],
			[f32(-0.128987), f32(0.70533),
				f32(0.685512)],
			[f32(-0.079877), f32(0.792123), f32(-0.591793)],
			[f32(-0.074164), f32(-0.867392),
				f32(-0.475594)],
			[f32(-0.001607), f32(0.156613), f32(0.979553)],
			[f32(0.001607), f32(-0.156613),
				f32(-0.979556)],
			[f32(0.074164), f32(0.867391), f32(0.475591)],
			[f32(0.079877), f32(-0.792124),
				f32(0.59179)],
			[f32(0.128987), f32(-0.70533), f32(-0.685515)],
			[f32(0.136047), f32(0.590601),
				f32(0.853427)],
			[f32(0.157929), f32(-0.433837), f32(-0.878011)],
			[f32(0.249306), f32(0.797226),
				f32(-0.535103)],
			[f32(0.255019), f32(-0.862289), f32(-0.418905)],
			[f32(0.280269), f32(-0.020452),
				f32(0.95136)],
			[f32(0.292369), f32(0.313377), f32(0.954971)],
			[f32(0.330629), f32(-0.606803),
				f32(0.711709)],
			[f32(0.33079), f32(-0.151511), f32(-0.922866)],
			[f32(0.339198), f32(0.752662),
				f32(0.643506)],
			[f32(0.373928), f32(0.858119), f32(0.328428)],
			[f32(0.37964), f32(-0.801396),
				f32(0.444627)],
			[f32(0.407172), f32(-0.312051), f32(0.849052)],
			[f32(0.482172), f32(0.814754),
				f32(-0.296215)],
			[f32(0.487884), f32(-0.844761), f32(-0.180016)],
			[f32(0.529773), f32(0.838013),
				f32(0.033625)],
			[f32(0.531183), f32(0.620161), f32(-0.563297)],
			[f32(0.535485), f32(-0.821502),
				f32(0.149823)],
			[f32(0.580033), f32(-0.029724), f32(0.804197)],
			[f32(0.581542), f32(0.03381),
				f32(-0.802948)],
			[f32(0.592133), f32(0.304105), f32(0.807809)],
			[f32(0.621074), f32(0.575598),
				f32(0.615313)],
			[f32(0.655804), f32(0.681055), f32(0.300235)],
			[f32(0.658086), f32(0.328562),
				f32(-0.665604)],
			[f32(0.738637), f32(-0.65944), f32(-0.060097)],
			[f32(0.783184), f32(0.132337),
				f32(0.594276)],
			[f32(0.812126), f32(0.40383), f32(0.40178)],
			[f32(0.814408), f32(0.051338), f32(-0.564059)],
			[f32(0.911497), f32(-0.377114),
				f32(-0.104953)],
			[f32(0.939029), f32(0.112232), f32(0.299472)],
			[f32(0.940439), f32(-0.10562),
				f32(-0.297449)],
			[f32(0.988041), f32(-0.082361), f32(0.032391)]]
		faces:    [[4, 8, 12], [3, 0, 1], [18, 28, 15], [9, 21, 16],
			[49, 45, 37], [52, 62, 55], [56, 43, 50], [64, 63, 67],
			[29, 23, 34], [36, 27, 31], [13, 19, 26], [5, 2, 6],
			[20, 32, 24], [7, 17, 14], [51, 54, 41], [60, 53, 48],
			[65, 57, 61], [69, 66, 68], [40, 35, 46], [33, 38, 42],
			[30, 40, 38], [22, 33, 21], [10, 9, 5], [13, 11, 6],
			[25, 26, 35], [58, 56, 63], [59, 64, 60], [47, 48, 36],
			[29, 39, 31], [44, 34, 43], [30, 25, 35, 40], [22, 30, 38, 33],
			[10, 22, 21, 9], [11, 10, 5, 6], [25, 11, 13, 26],
			[58, 44, 43, 56], [59, 58, 63, 64], [47, 59, 60, 48],
			[39, 47, 36, 31], [44, 39, 29, 34], [25, 30, 22, 10, 11],
			[44, 58, 59, 47, 39], [15, 28, 37, 45, 50, 43, 34, 23, 12, 8],
			[5, 9, 16, 18, 15, 8, 4, 1, 0, 2], [42, 52, 55, 49, 37, 28, 18, 16, 21, 33],
			[69, 67, 63, 56, 50, 45, 49, 55, 62, 66], [67, 69, 68, 65, 61, 54, 51, 53, 60, 64],
			[7, 3, 1, 4, 12, 23, 29, 31, 27, 17], [24, 32, 41, 54, 61, 57, 46, 35, 26, 19],
			[3, 7, 14, 20, 24, 19, 13, 6, 2, 0], [36, 48, 53, 51, 41, 32, 20, 14, 17, 27],
			[52, 42, 38, 40, 46, 57, 65, 68, 66, 62]]
	},
	&Polyhedron{
		name:     'j70'
		vertexes: [[f32(-0.989194), f32(-0.091477), f32(-0.102373)],
			[f32(-0.986156), f32(-0.109996), f32(0.232129)],
			[f32(-0.908902), f32(0.23333),
				f32(-0.08512)],
			[f32(-0.905864), f32(0.214811), f32(0.249382)],
			[f32(-0.892465), f32(-0.388533),
				f32(-0.22339)],
			[f32(-0.887549), f32(-0.418497), f32(0.317846)],
			[f32(-0.850998), f32(0.061184),
				f32(-0.366646)],
			[f32(-0.843044), f32(0.012701), f32(0.509091)],
			[f32(-0.829645), f32(-0.590642),
				f32(0.03632)],
			[f32(-0.810408), f32(0.497156), f32(0.096369)],
			[f32(-0.754269), f32(-0.235871),
				f32(-0.487662)],
			[f32(-0.744438), f32(-0.2958), f32(0.594808)],
			[f32(-0.658813), f32(0.046474),
				f32(-0.640675)],
			[f32(-0.655662), f32(-0.544372), f32(-0.401946)],
			[f32(-0.647709), f32(-0.592856), f32(0.473792)],
			[f32(-0.645943), f32(-0.031974),
				f32(0.776297)],
			[f32(-0.593136), f32(0.75189), f32(0.108498)],
			[f32(-0.592842), f32(-0.746482),
				f32(-0.142236)],
			[f32(-0.589804), f32(-0.765001), f32(0.192266)],
			[f32(-0.405755), f32(0.194817),
				f32(-0.802538)],
			[f32(-0.400657), f32(-0.761193), f32(-0.416265)],
			[f32(-0.392703), f32(-0.809676), f32(0.459472)],
			[f32(-0.389847), f32(0.09785),
				f32(0.948936)],
			[f32(-0.340078), f32(0.900233), f32(-0.053365)],
			[f32(-0.33704), f32(0.881715),
				f32(0.281137)],
			[f32(-0.188483), f32(0.449551), f32(-0.790409)],
			[f32(-0.172576), f32(0.352585),
				f32(0.961066)],
			[f32(-0.147893), f32(0.885523), f32(-0.327394)],
			[f32(-0.139939), f32(0.83704),
				f32(0.548343)],
			[f32(-0.091754), f32(0.152496), f32(-0.911425)],
			[f32(-0.089989), f32(0.713378),
				f32(-0.60892)],
			[f32(-0.086657), f32(-0.803514), f32(-0.525152)],
			[f32(-0.07712), f32(0.63493), f32(0.808053)],
			[f32(-0.076826), f32(-0.863443),
				f32(0.557318)],
			[f32(-0.073969), f32(0.044084), f32(1.04678)],
			[f32(0.126005), f32(0.562254),
				f32(-0.815685)],
			[f32(0.163251), f32(-0.064325), f32(-0.925745)],
			[f32(0.166107), f32(0.843202),
				f32(-0.436281)],
			[f32(0.166401), f32(-0.655171), f32(-0.687015)],
			[f32(0.175938), f32(0.783273),
				f32(0.64619)],
			[f32(0.179271), f32(-0.733618), f32(0.729957)],
			[f32(0.181036), f32(-0.172737),
				f32(1.03246)],
			[f32(0.222734), f32(0.265199), f32(-0.936702)],
			[f32(0.229221), f32(-0.857281),
				f32(-0.427306)],
			[f32(0.237175), f32(-0.905764), f32(0.448431)],
			[f32(0.261857), f32(-0.372826),
				f32(-0.840028)],
			[f32(0.277765), f32(-0.469792), f32(0.911446)],
			[f32(0.382101), f32(0.692078),
				f32(-0.643046)],
			[f32(0.426322), f32(-0.901955), f32(-0.1601)],
			[f32(0.42936), f32(-0.920474),
				f32(0.174402)],
			[f32(0.479129), f32(-0.118091), f32(-0.827899)],
			[f32(0.481985), f32(0.789435),
				f32(-0.338434)],
			[f32(0.489939), f32(0.740952), f32(0.537303)],
			[f32(0.495036), f32(-0.215058),
				f32(0.923576)],
			[f32(0.538612), f32(0.211432), f32(-0.838855)],
			[f32(0.637106), f32(0.475258),
				f32(-0.657366)],
			[f32(0.679086), f32(0.74476), f32(-0.071228)],
			[f32(0.682124), f32(0.726241),
				f32(0.263273)],
			[f32(0.682418), f32(-0.772131), f32(0.012539)],
			[f32(0.735225), f32(0.011733),
				f32(-0.65526)],
			[f32(0.73699), f32(0.572615), f32(-0.352754)],
			[f32(0.744944), f32(0.524132),
				f32(0.522983)],
			[f32(0.748094), f32(-0.066715), f32(0.761713)],
			[f32(0.833719), f32(0.275559),
				f32(-0.473771)],
			[f32(0.84355), f32(0.21563), f32(0.6087)], [f32(0.899689), f32(-0.517397), f32(0.024669)],
			[f32(0.932326), f32(-0.032942), f32(-0.388054)],
			[f32(0.940279), f32(-0.081425),
				f32(0.487683)],
			[f32(0.995146), f32(-0.235051), f32(-0.128344)],
			[f32(0.998184), f32(-0.253571),
				f32(0.206158)]]
		faces:    [[41, 46, 53], [26, 22, 34], [33, 44, 40], [14, 18, 21],
			[48, 58, 49], [31, 38, 43], [68, 69, 65], [59, 63, 66],
			[64, 62, 67], [57, 52, 61], [3, 9, 2], [11, 15, 7],
			[24, 23, 16], [32, 39, 28], [37, 30, 27], [60, 51, 56],
			[29, 19, 25], [50, 45, 36], [10, 6, 12], [17, 13, 20],
			[4, 10, 13], [8, 17, 18], [5, 14, 11], [3, 1, 7],
			[0, 2, 6], [47, 37, 51], [55, 60, 63], [54, 59, 50],
			[29, 42, 36], [35, 25, 30], [4, 0, 6, 10], [8, 4, 13, 17],
			[5, 8, 18, 14], [1, 5, 11, 7], [0, 1, 3, 2], [47, 35, 30, 37],
			[55, 47, 51, 60], [54, 55, 63, 59], [42, 54, 50, 36],
			[35, 42, 29, 25], [0, 4, 8, 5, 1], [35, 47, 55, 54, 42],
			[40, 44, 49, 58, 65, 69, 67, 62, 53, 46], [11, 14, 21, 33, 40, 46, 41, 34, 22, 15],
			[20, 31, 43, 48, 49, 44, 33, 21, 18, 17], [50, 59, 66, 68, 65, 58, 48, 43, 38, 45],
			[56, 57, 61, 64, 67, 69, 68, 66, 63, 60], [32, 26, 34, 41, 53, 62, 64, 61, 52, 39],
			[16, 23, 27, 30, 25, 19, 12, 6, 2, 9], [26, 32, 28, 24, 16, 9, 3, 7, 15, 22],
			[57, 56, 51, 37, 27, 23, 24, 28, 39, 52], [31, 20, 13, 10, 12, 19, 29, 36, 45, 38]]
	},
	&Polyhedron{
		name:     'j71'
		vertexes: [[f32(-0.942902), f32(0.07027), f32(-0.149675)],
			[f32(-0.907058), f32(0.322313), f32(0.065363)],
			[f32(-0.897048), f32(-0.257164),
				f32(-0.191336)],
			[f32(-0.851819), f32(0.371393), f32(-0.259585)],
			[f32(-0.803207), f32(0.402693),
				f32(0.37164)],
			[f32(-0.802539), f32(0.632087), f32(0.129919)],
			[f32(-0.787011), f32(-0.534922),
				f32(-0.043707)],
			[f32(-0.7473), f32(0.681167), f32(-0.195029)],
			[f32(-0.731772), f32(-0.485841),
				f32(-0.368655)],
			[f32(-0.671018), f32(0.280706), f32(0.65217)],
			[f32(-0.658589), f32(0.531186),
				f32(-0.479085)],
			[f32(-0.654821), f32(-0.656908), f32(0.236823)],
			[f32(-0.579935), f32(0.581829),
				f32(0.542259)],
			[f32(-0.579266), f32(0.811224), f32(0.300537)],
			[f32(-0.560981), f32(0.002949),
				f32(0.799799)],
			[f32(-0.550971), f32(-0.576528), f32(0.5431)],
			[f32(-0.515127), f32(-0.324486),
				f32(0.758138)],
			[f32(-0.510203), f32(-0.528414), f32(-0.613902)],
			[f32(-0.489887), f32(0.890637), f32(-0.225239)],
			[f32(-0.437021), f32(0.488613),
				f32(-0.724333)],
			[f32(-0.401177), f32(0.740656), f32(-0.509295)],
			[f32(-0.386037), f32(0.971017),
				f32(0.081037)],
			[f32(-0.385694), f32(-0.805205), f32(0.365781)],
			[f32(-0.322522), f32(0.791299),
				f32(0.512049)],
			[f32(-0.317618), f32(-0.591958), f32(0.780503)],
			[f32(-0.316974), f32(-0.368621),
				f32(-0.833402)],
			[f32(-0.291854), f32(-0.145349), f32(0.928756)],
			[f32(-0.271745), f32(0.259936),
				f32(-0.901652)],
			[f32(-0.225891), f32(-0.067498), f32(-0.943313)],
			[f32(-0.206937), f32(-0.646378), f32(-0.685774)],
			[f32(-0.177904), f32(0.919793), f32(-0.338677)],
			[f32(-0.152342), f32(-0.820635),
				f32(0.603184)],
			[f32(-0.129293), f32(0.951092), f32(0.292549)],
			[f32(-0.094345), f32(-0.412822),
				f32(0.951122)],
			[f32(-0.082428), f32(-0.92317), f32(0.29391)],
			[f32(-0.074054), f32(1.00017),
				f32(-0.032399)],
			[f32(0.002897), f32(0.829106), f32(0.573078)],
			[f32(0.031522), f32(0.141972),
				f32(-0.973523)],
			[f32(0.033565), f32(-0.107542), f32(0.989786)],
			[f32(0.06219), f32(-0.794676),
				f32(-0.556816)],
			[f32(0.13914), f32(-0.965743), f32(0.048662)],
			[f32(0.147515), f32(0.9576), f32(-0.277647)],
			[f32(0.173077), f32(-0.782829),
				f32(0.664213)],
			[f32(0.19438), f32(-0.916662), f32(-0.276286)],
			[f32(0.208921), f32(-0.530786),
				f32(0.87925)],
			[f32(0.242991), f32(-0.885363), f32(0.354939)],
			[f32(0.272024), f32(0.680808),
				f32(0.702036)],
			[f32(0.290978), f32(0.101928), f32(0.959576)],
			[f32(0.336832), f32(-0.225507),
				f32(0.917915)],
			[f32(0.356941), f32(0.179778), f32(-0.912493)],
			[f32(0.382061), f32(0.403051),
				f32(0.849665)],
			[f32(0.387609), f32(-0.75687), f32(-0.495786)],
			[f32(0.450781), f32(0.839635),
				f32(-0.349518)],
			[f32(0.466264), f32(-0.706226), f32(0.525558)],
			[f32(0.502108), f32(-0.454184),
				f32(0.740596)],
			[f32(0.57529), f32(0.562844), f32(0.630165)],
			[f32(0.580214), f32(0.358915),
				f32(-0.741875)],
			[f32(-0.018946), f32(-0.326587), f32(-0.976456)],
			[f32(0.616058), f32(0.610958), f32(-0.526838)],
			[f32(0.626068), f32(0.031481),
				f32(-0.783536)],
			[f32(0.645022), f32(-0.5474), f32(-0.525996)],
			[f32(0.238466), f32(-0.117117),
				f32(-1.00667)],
			[f32(0.719908), f32(0.691337), f32(-0.22056)],
			[f32(0.723676), f32(-0.496756),
				f32(0.495348)],
			[f32(0.736105), f32(-0.246276), f32(-0.635907)],
			[f32(0.796859), f32(0.520271),
				f32(0.384917)],
			[f32(0.091091), f32(-0.604344), f32(-0.828827)],
			[f32(0.852098), f32(0.569351),
				f32(0.059969)],
			[f32(0.868294), f32(-0.368263), f32(-0.355377)],
			[f32(0.507593), f32(-0.265415),
				f32(-0.877708)],
			[f32(0.916906), f32(-0.336964), f32(0.275848)],
			[f32(0.962135), f32(0.291594),
				f32(0.207599)],
			[f32(0.41651), f32(-0.566538), f32(-0.767798)],
			[f32(0.972145), f32(-0.287883),
				f32(-0.0491)],
			[f32(1.00799), f32(-0.035841), f32(0.165937)]]
		faces:    [[70, 73, 74], [54, 53, 63], [60, 64, 68], [43, 39, 51],
			[49, 56, 59], [28, 27, 37], [52, 62, 58], [30, 35, 41],
			[65, 71, 67], [50, 55, 46], [3, 0, 1], [20, 19, 10],
			[8, 6, 2], [25, 29, 17], [22, 15, 11], [45, 34, 40],
			[26, 14, 16], [48, 47, 38], [12, 4, 9], [32, 23, 36],
			[13, 12, 23], [21, 32, 35], [18, 30, 20], [3, 7, 10],
			[5, 1, 4], [31, 22, 34], [42, 45, 53], [44, 54, 48],
			[26, 33, 38], [24, 16, 15], [66, 39, 29], [57, 25, 28],
			[61, 37, 49], [69, 59, 64], [72, 60, 51], [13, 5, 4, 12],
			[21, 13, 23, 32], [18, 21, 35, 30], [7, 18, 20, 10],
			[5, 7, 3, 1], [31, 24, 15, 22], [42, 31, 34, 45],
			[44, 42, 53, 54], [33, 44, 48, 38], [24, 33, 26, 16],
			[66, 72, 51, 39], [66, 29, 25, 57], [57, 28, 37, 61],
			[61, 49, 59, 69], [69, 64, 60, 72], [5, 13, 21, 18, 7],
			[24, 31, 42, 44, 33], [72, 66, 57, 61, 69], [68, 64, 59, 56, 58, 62, 67, 71, 74, 73],
			[40, 43, 51, 60, 68, 73, 70, 63, 53, 45], [54, 63, 70, 74, 71, 65, 55, 50, 47, 48],
			[20, 30, 41, 52, 58, 56, 49, 37, 27, 19], [36, 46, 55, 65, 67, 62, 52, 41, 35, 32],
			[2, 6, 11, 15, 16, 14, 9, 4, 1, 0], [28, 25, 17, 8, 2, 0, 3, 10, 19, 27],
			[43, 40, 34, 22, 11, 6, 8, 17, 29, 39], [46, 36, 23, 12, 9, 14, 26, 38, 47, 50]]
	},
	&Polyhedron{
		name:     'j72'
		vertexes: [[f32(-0.976612), f32(0.213547), f32(-0.025026)],
			[f32(-0.942883), f32(-0.134569), f32(-0.304734)],
			[f32(-0.917763), f32(0.061996), f32(0.392261)],
			[f32(-0.863187), f32(-0.501268),
				f32(-0.060316)],
			[f32(-0.847662), f32(-0.379783), f32(0.37045)],
			[f32(-0.806942), f32(0.483006),
				f32(-0.339927)],
			[f32(-0.791417), f32(0.60449), f32(0.090839)],
			[f32(-0.773213), f32(0.13489),
				f32(-0.619635)],
			[f32(-0.732567), f32(0.452939), f32(0.508126)],
			[f32(-0.703113), f32(-0.306889),
				f32(-0.641445)],
			[f32(-0.652871), f32(0.086241), f32(0.752543)],
			[f32(-0.623417), f32(-0.673588),
				f32(-0.397028)],
			[f32(-0.582771), f32(-0.355538), f32(0.730732)],
			[f32(-0.564567), f32(-0.825138),
				f32(0.020258)],
			[f32(-0.549042), f32(-0.703654), f32(0.451025)],
			[f32(-0.47356), f32(0.76745),
				f32(-0.432161)],
			[f32(-0.458035), f32(0.888934), f32(-0.001394)],
			[f32(-0.418985), f32(0.204186),
				f32(-0.884738)],
			[f32(-0.362814), f32(0.643719), f32(0.673789)],
			[f32(-0.348885), f32(-0.237593),
				f32(-0.906548)],
			[f32(-0.283118), f32(0.277021), f32(0.918206)],
			[f32(-0.23379), f32(0.595129),
				f32(-0.768872)],
			[f32(-0.219935), f32(-0.830923), f32(-0.511073)],
			[f32(-0.193143), f32(0.913179), f32(0.358888)],
			[f32(-0.169693), f32(-0.437793),
				f32(0.882916)],
			[f32(-0.161085), f32(-0.982474), f32(-0.093786)],
			[f32(-0.135964), f32(-0.785909), f32(0.603208)],
			[f32(-0.103807), f32(0.95823),
				f32(-0.266497)],
			[f32(-0.050264), f32(-0.561464), f32(-0.825973)],
			[f32(-0.015503), f32(0.04685), f32(-0.998782)],
			[f32(0.015502), f32(-0.04685),
				f32(0.998781)],
			[f32(0.075132), f32(0.737294), f32(0.671381)],
			[f32(0.103807), f32(-0.958229),
				f32(0.266497)],
			[f32(0.135964), f32(0.78591), f32(-0.603209)],
			[f32(0.154828), f32(0.370596),
				f32(0.915798)],
			[f32(0.161084), f32(0.982475), f32(0.093785)],
			[f32(0.169693), f32(0.437794),
				f32(-0.882917)],
			[f32(0.193143), f32(-0.913178), f32(-0.358889)],
			[f32(0.233789), f32(-0.595129),
				f32(0.768871)],
			[f32(0.283118), f32(-0.277021), f32(-0.918207)],
			[f32(0.362813), f32(-0.643719),
				f32(-0.67379)],
			[f32(0.418985), f32(-0.204186), f32(0.884737)],
			[f32(0.42936), f32(0.80659), f32(0.406278)],
			[f32(0.458035), f32(-0.888933), f32(0.001394)],
			[f32(0.47356), f32(-0.767449),
				f32(0.43216)],
			[f32(0.549042), f32(0.703655), f32(-0.451025)],
			[f32(0.558311), f32(0.21326),
				f32(0.801754)],
			[f32(0.564567), f32(0.825139), f32(-0.020259)],
			[f32(0.582771), f32(0.355539),
				f32(-0.730733)],
			[f32(0.652871), f32(-0.08624), f32(-0.752544)],
			[f32(0.727981), f32(0.48272),
				f32(0.486853)],
			[f32(0.732567), f32(-0.452939), f32(-0.508127)],
			[f32(0.773213), f32(-0.13489),
				f32(0.619634)],
			[f32(0.791417), f32(-0.60449), f32(-0.09084)],
			[f32(0.806942), f32(-0.483006),
				f32(0.339926)],
			[f32(0.847662), f32(0.379784), f32(-0.370451)],
			[f32(0.863187), f32(0.501268),
				f32(0.060316)],
			[f32(0.917763), f32(-0.061995), f32(-0.392261)],
			[f32(0.942883), f32(0.13457),
				f32(0.304733)],
			[f32(0.976612), f32(-0.213546), f32(0.025025)]]
		faces:    [[48, 45, 55], [35, 42, 47], [23, 18, 31], [20, 30, 34],
			[49, 57, 51], [59, 54, 53], [56, 50, 58], [46, 41, 52],
			[39, 40, 28], [37, 25, 22], [43, 44, 32], [38, 24, 26],
			[29, 19, 17], [9, 1, 7], [11, 13, 3], [14, 12, 4],
			[36, 21, 33], [15, 16, 27], [5, 0, 6], [2, 10, 8],
			[36, 33, 45, 48], [45, 47, 56, 55], [47, 42, 50, 56],
			[23, 31, 42, 35], [18, 20, 34, 31], [34, 30, 41, 46],
			[48, 55, 57, 49], [57, 59, 53, 51], [53, 54, 44, 43],
			[58, 52, 54, 59], [50, 46, 52, 58], [41, 30, 24, 38],
			[49, 51, 40, 39], [40, 37, 22, 28], [22, 25, 13, 11],
			[43, 32, 25, 37], [44, 38, 26, 32], [26, 24, 12, 14],
			[39, 28, 19, 29], [19, 9, 7, 17], [7, 1, 0, 5], [11, 3, 1, 9],
			[13, 14, 4, 3], [4, 12, 10, 2], [29, 17, 21, 36],
			[21, 15, 27, 33], [27, 16, 23, 35], [5, 6, 16, 15],
			[0, 2, 8, 6], [8, 10, 20, 18], [33, 27, 35, 47, 45],
			[31, 34, 46, 50, 42], [55, 56, 58, 59, 57], [52, 41, 38, 44, 54],
			[51, 53, 43, 37, 40], [32, 26, 14, 13, 25], [28, 22, 11, 9, 19],
			[3, 4, 2, 0, 1], [17, 7, 5, 15, 21], [6, 8, 18, 23, 16],
			[36, 48, 49, 39, 29], [10, 12, 24, 30, 20]]
	},
	&Polyhedron{
		name:     'j73'
		vertexes: [[f32(-0.984691), f32(0.125192), f32(0.121281)],
			[f32(-0.957572), f32(-0.075612), f32(-0.278094)],
			[f32(-0.942455), f32(-0.319982), f32(0.096891)],
			[f32(-0.856557), f32(0.512005),
				f32(-0.064506)],
			[f32(-0.832097), f32(0.116607), f32(0.542233)],
			[f32(-0.829438), f32(0.3112),
				f32(-0.463882)],
			[f32(-0.789861), f32(-0.328568), f32(0.517842)],
			[f32(-0.761099), f32(-0.409107),
				f32(-0.503346)],
			[f32(-0.745982), f32(-0.653477), f32(-0.128361)],
			[f32(-0.624772), f32(0.742482), f32(0.241623)],
			[f32(-0.609655), f32(0.498112),
				f32(0.616608)],
			[f32(-0.606996), f32(0.692705), f32(-0.389506)],
			[f32(-0.558076), f32(-0.098091),
				f32(0.823971)],
			[f32(-0.553774), f32(0.216768), f32(-0.803956)],
			[f32(-0.511538), f32(-0.228406),
				f32(-0.828346)],
			[f32(-0.49908), f32(-0.667369), f32(0.552753)],
			[f32(-0.471962), f32(-0.868174),
				f32(0.153378)],
			[f32(-0.40552), f32(-0.630422), f32(-0.661906)],
			[f32(-0.390403), f32(-0.874792),
				f32(-0.286921)],
			[f32(-0.375211), f32(0.923183), f32(-0.083378)],
			[f32(-0.335634), f32(0.283415),
				f32(0.898346)],
			[f32(-0.331332), f32(0.598273), f32(-0.729581)],
			[f32(-0.287416), f32(0.79711),
				f32(0.531045)],
			[f32(-0.267295), f32(-0.436892), f32(0.858882)],
			[f32(-0.134858), f32(0.264778),
				f32(-0.954832)],
			[f32(-0.092623), f32(-0.180396), f32(-0.979223)],
			[f32(-0.070822), f32(-0.770387), f32(0.63363)],
			[f32(-0.043703), f32(-0.971192),
				f32(0.234255)],
			[f32(-0.037854), f32(0.977811), f32(0.206045)],
			[f32(-0.013394), f32(0.582413),
				f32(0.812784)],
			[f32(0.013396), f32(-0.582411), f32(-0.812783)],
			[f32(0.037856), f32(-0.977809),
				f32(-0.206044)],
			[f32(0.043705), f32(0.971193), f32(-0.234254)],
			[f32(0.070824), f32(0.770388),
				f32(-0.63363)],
			[f32(0.092624), f32(0.180397), f32(0.979223)],
			[f32(0.13486), f32(-0.264777),
				f32(0.954833)],
			[f32(0.267297), f32(0.436893), f32(-0.858881)],
			[f32(0.287417), f32(-0.797109),
				f32(-0.531044)],
			[f32(0.331333), f32(-0.598272), f32(0.729581)],
			[f32(0.335635), f32(-0.283414),
				f32(-0.898346)],
			[f32(0.375212), f32(-0.923181), f32(0.083378)],
			[f32(0.390404), f32(0.874793),
				f32(0.286922)],
			[f32(0.405521), f32(0.630423), f32(0.661907)],
			[f32(0.471963), f32(0.868175),
				f32(-0.153377)],
			[f32(0.499082), f32(0.66737), f32(-0.552753)],
			[f32(0.511539), f32(0.228408),
				f32(0.828347)],
			[f32(0.553775), f32(-0.216766), f32(0.803957)],
			[f32(0.558078), f32(0.098092),
				f32(-0.823971)],
			[f32(0.606997), f32(-0.692704), f32(0.389507)],
			[f32(0.609656), f32(-0.498111),
				f32(-0.616607)],
			[f32(0.624773), f32(-0.74248), f32(-0.241622)],
			[f32(0.745984), f32(0.653478),
				f32(0.128361)],
			[f32(0.761101), f32(0.409108), f32(0.503346)],
			[f32(0.789863), f32(0.328569),
				f32(-0.517842)],
			[f32(0.82944), f32(-0.311199), f32(0.463882)],
			[f32(0.832099), f32(-0.116605),
				f32(-0.542232)],
			[f32(0.856558), f32(-0.512003), f32(0.064507)],
			[f32(0.942457), f32(0.319983),
				f32(-0.09689)],
			[f32(0.957574), f32(0.075614), f32(0.278095)],
			[f32(0.984692), f32(-0.125191),
				f32(-0.121281)]]
		faces:    [[36, 33, 44], [19, 28, 32], [9, 10, 22], [20, 34, 29],
			[47, 53, 55], [57, 58, 59], [43, 41, 51], [42, 45, 52],
			[49, 50, 37], [40, 27, 31], [56, 54, 48], [46, 35, 38],
			[39, 30, 25], [17, 7, 14], [18, 16, 8], [26, 23, 15],
			[24, 13, 21], [5, 3, 11], [1, 2, 0], [6, 12, 4], [24, 21, 33, 36],
			[33, 32, 43, 44], [32, 28, 41, 43], [9, 22, 28, 19],
			[10, 20, 29, 22], [29, 34, 45, 42], [36, 44, 53, 47],
			[53, 57, 59, 55], [59, 58, 54, 56], [51, 52, 58, 57],
			[41, 42, 52, 51], [45, 34, 35, 46], [47, 55, 49, 39],
			[50, 40, 31, 37], [31, 27, 16, 18], [56, 48, 40, 50],
			[54, 46, 38, 48], [38, 35, 23, 26], [49, 37, 30, 39],
			[30, 17, 14, 25], [7, 8, 2, 1], [18, 8, 7, 17], [27, 26, 15, 16],
			[15, 23, 12, 6], [25, 14, 13, 24], [13, 5, 11, 21],
			[11, 3, 9, 19], [1, 0, 3, 5], [2, 6, 4, 0], [4, 12, 20, 10],
			[21, 11, 19, 32, 33], [22, 29, 42, 41, 28], [44, 43, 51, 57, 53],
			[52, 45, 46, 54, 58], [55, 59, 56, 50, 49], [48, 38, 26, 27, 40],
			[37, 31, 18, 17, 30], [16, 15, 6, 2, 8], [14, 7, 1, 5, 13],
			[0, 4, 10, 9, 3], [24, 36, 47, 39, 25], [12, 23, 35, 34, 20]]
	},
	&Polyhedron{
		name:     'j74'
		vertexes: [[f32(-0.966046), f32(-0.051368), f32(0.253213)],
			[f32(-0.95229), f32(0.30466), f32(-0.018105)],
			[f32(-0.940892), f32(-0.323),
				f32(-0.101952)],
			[f32(-0.927135), f32(0.033028), f32(-0.37327)],
			[f32(-0.826492), f32(-0.473879),
				f32(0.30389)],
			[f32(-0.790478), f32(0.458215), f32(-0.40643)],
			[f32(-0.767188), f32(0.060532),
				f32(0.63856)],
			[f32(-0.744929), f32(0.636598), f32(0.199559)],
			[f32(-0.701332), f32(-0.650609),
				f32(-0.291274)],
			[f32(-0.679074), f32(-0.074543), f32(-0.730275)],
			[f32(-0.63053), f32(0.485719), f32(0.6054)],
			[f32(-0.627634), f32(-0.361979),
				f32(0.689237)],
			[f32(-0.586933), f32(-0.801488), f32(0.114568)],
			[f32(-0.583117), f32(0.790154),
				f32(-0.188766)],
			[f32(-0.542416), f32(0.350644), f32(-0.763435)],
			[f32(-0.53952), f32(-0.497054),
				f32(-0.679599)],
			[f32(-0.420274), f32(-0.03004), f32(0.9069)],
			[f32(-0.397364), f32(0.817911),
				f32(0.416083)],
			[f32(-0.338872), f32(-0.909059), f32(-0.242438)],
			[f32(-0.302857), f32(0.023036), f32(-0.952757)],
			[f32(-0.283617), f32(0.395147),
				f32(0.87374)],
			[f32(-0.265174), f32(-0.620429), f32(0.738072)],
			[f32(-0.240019), f32(-0.892061),
				f32(0.382907)],
			[f32(-0.235552), f32(0.971466), f32(0.027758)],
			[f32(-0.206901), f32(0.887732),
				f32(-0.411248)],
			[f32(-0.181746), f32(0.6161), f32(-0.766413)],
			[f32(-0.17706), f32(-0.755504),
				f32(-0.630763)],
			[f32(-0.163303), f32(-0.399475), f32(-0.902081)],
			[f32(-0.057814), f32(-0.288491), f32(0.955736)],
			[f32(-0.05045), f32(0.727338),
				f32(0.684423)],
			[f32(0.008042), f32(-0.999632), f32(0.025902)],
			[f32(0.057813), f32(0.288491),
				f32(-0.955736)],
			[f32(0.163303), f32(0.399477), f32(0.902082)],
			[f32(0.181745), f32(-0.616099),
				f32(0.766414)],
			[f32(0.2069), f32(-0.887731), f32(0.411249)], [f32(0.211368), f32(0.975796), f32(0.0561)],
			[f32(0.240019), f32(0.892062), f32(-0.382907)],
			[f32(0.265173), f32(0.62043),
				f32(-0.738072)],
			[f32(0.26986), f32(-0.751174), f32(-0.602422)],
			[f32(0.283616), f32(-0.395146),
				f32(-0.873739)],
			[f32(0.302857), f32(-0.023034), f32(0.952758)],
			[f32(0.325767), f32(0.824917),
				f32(0.461941)],
			[f32(0.384259), f32(-0.902053), f32(-0.19658)],
			[f32(0.420273), f32(0.030041),
				f32(-0.9069)],
			[f32(0.539519), f32(0.497055), f32(0.6796)],
			[f32(0.542416), f32(-0.350643), f32(0.763436)],
			[f32(0.583117), f32(-0.790152),
				f32(0.188767)],
			[f32(0.586933), f32(0.801489), f32(-0.114567)],
			[f32(0.627634), f32(0.36198),
				f32(-0.689236)],
			[f32(0.658347), f32(-0.625824), f32(-0.418238)],
			[f32(0.672103), f32(-0.269795),
				f32(-0.689555)],
			[f32(0.679073), f32(0.074544), f32(0.730276)],
			[f32(0.701332), f32(0.65061), f32(0.291275)],
			[f32(0.790477), f32(-0.458214), f32(0.40643)],
			[f32(0.826492), f32(0.473881),
				f32(-0.303889)],
			[f32(0.857205), f32(-0.513923), f32(-0.03289)],
			[f32(0.879463), f32(0.062143),
				f32(-0.471892)],
			[f32(0.927134), f32(-0.033027), f32(0.37327)],
			[f32(0.940891), f32(0.323002),
				f32(0.101953)],
			[f32(0.993863), f32(-0.088736), f32(-0.06605)]]
		faces:    [[31, 25, 37], [13, 23, 24], [7, 10, 17], [20, 32, 29],
			[48, 54, 56], [58, 57, 59], [36, 35, 47], [41, 44, 52],
			[43, 50, 39], [49, 42, 38], [55, 53, 46], [51, 40, 45],
			[27, 26, 15], [18, 12, 8], [30, 34, 22], [33, 28, 21],
			[19, 9, 14], [3, 1, 5], [2, 4, 0], [11, 16, 6], [19, 14, 25, 31],
			[25, 24, 36, 37], [24, 23, 35, 36], [7, 17, 23, 13],
			[10, 20, 29, 17], [29, 32, 44, 41], [31, 37, 48, 43],
			[54, 58, 59, 56], [59, 57, 53, 55], [47, 52, 58, 54],
			[35, 41, 52, 47], [44, 32, 40, 51], [48, 56, 50, 43],
			[50, 49, 38, 39], [42, 46, 34, 30], [55, 46, 42, 49],
			[57, 51, 45, 53], [45, 40, 28, 33], [39, 38, 26, 27],
			[26, 18, 8, 15], [8, 12, 4, 2], [30, 22, 12, 18],
			[34, 33, 21, 22], [21, 28, 16, 11], [27, 15, 9, 19],
			[9, 3, 5, 14], [5, 1, 7, 13], [2, 0, 1, 3], [4, 11, 6, 0],
			[6, 16, 20, 10], [14, 5, 13, 24, 25], [17, 29, 41, 35, 23],
			[37, 36, 47, 54, 48], [52, 44, 51, 57, 58], [56, 59, 55, 49, 50],
			[53, 45, 33, 34, 46], [38, 42, 30, 18, 26], [22, 21, 11, 4, 12],
			[15, 8, 2, 3, 9], [0, 6, 10, 7, 1], [19, 31, 43, 39, 27],
			[16, 28, 40, 32, 20]]
	},
	&Polyhedron{
		name:     'j75'
		vertexes: [[f32(-0.980376), f32(-0.197048), f32(-0.005857)],
			[f32(-0.946332), f32(0.150802), f32(-0.285858)],
			[f32(-0.935804), f32(0.079716),
				f32(0.34339)],
			[f32(-0.901759), f32(0.427566), f32(0.063389)],
			[f32(-0.812124), f32(-0.53251),
				f32(0.23851)],
			[f32(-0.8048), f32(-0.555655), f32(-0.20867)],
			[f32(-0.767552), f32(-0.255746),
				f32(0.587757)],
			[f32(-0.759203), f32(0.553784), f32(-0.341957)],
			[f32(-0.749715), f32(0.007177),
				f32(-0.661721)],
			[f32(-0.688108), f32(0.168923), f32(0.705672)],
			[f32(-0.662244), f32(-0.429437),
				f32(-0.614016)],
			[f32(-0.633023), f32(0.731755), f32(0.252621)],
			[f32(-0.562586), f32(0.41016),
				f32(-0.71782)],
			[f32(-0.500979), f32(0.571905), f32(0.649573)],
			[f32(-0.490467), f32(0.857973),
				f32(-0.152725)],
			[f32(-0.483464), f32(-0.835984), f32(0.259599)],
			[f32(-0.47614), f32(-0.859129),
				f32(-0.18758)],
			[f32(-0.411344), f32(-0.388171), f32(0.824694)],
			[f32(-0.387011), f32(0.051553),
				f32(-0.920632)],
			[f32(-0.333584), f32(-0.732911), f32(-0.592926)],
			[f32(-0.331901), f32(0.036498), f32(0.942608)],
			[f32(-0.299539), f32(-0.385062),
				f32(-0.872928)],
			[f32(-0.245677), f32(0.868112), f32(0.431306)],
			[f32(-0.235768), f32(-0.746778),
				f32(0.621881)],
			[f32(-0.172335), f32(0.625585), f32(-0.760884)],
			[f32(-0.144772), f32(0.43948),
				f32(0.88651)],
			[f32(-0.127762), f32(0.902348), f32(-0.411637)],
			[f32(-0.119933), f32(-0.991554),
				f32(0.049356)],
			[f32(-0.103121), f32(0.994331), f32(0.02596)],
			[f32(-0.003241), f32(-0.266976),
				f32(0.963698)],
			[f32(0.003241), f32(0.266978), f32(-0.963697)],
			[f32(0.11053), f32(0.735688),
				f32(0.668243)],
			[f32(0.110728), f32(-0.787329), f32(-0.606508)],
			[f32(0.127763), f32(-0.902347),
				f32(0.411638)],
			[f32(0.144773), f32(-0.439479), f32(-0.886509)],
			[f32(0.172335), f32(-0.625583),
				f32(0.760885)],
			[f32(0.242772), f32(-0.947178), f32(-0.209555)],
			[f32(0.271977), f32(0.571167),
				f32(-0.774465)],
			[f32(0.29954), f32(0.385063), f32(0.872928)],
			[f32(0.31655), f32(0.847931), f32(-0.425218)],
			[f32(0.331901), f32(-0.036497),
				f32(-0.942608)],
			[f32(0.341191), f32(0.939913), f32(0.012379)],
			[f32(0.387011), f32(-0.051552),
				f32(0.920633)],
			[f32(0.473235), f32(0.780063), f32(0.409331)],
			[f32(0.490467), f32(-0.857972),
				f32(0.152726)],
			[f32(0.528066), f32(-0.712229), f32(-0.462467)],
			[f32(0.562111), f32(-0.364379),
				f32(-0.742468)],
			[f32(0.562587), f32(-0.410159), f32(0.717821)],
			[f32(0.600637), f32(0.267692),
				f32(-0.753376)],
			[f32(0.662244), f32(0.429438), f32(0.614017)],
			[f32(0.672757), f32(0.715506),
				f32(-0.188282)],
			[f32(0.749716), f32(-0.007176), f32(0.661722)],
			[f32(0.759203), f32(-0.553783),
				f32(0.341958)],
			[f32(0.775762), f32(-0.623022), f32(-0.100185)],
			[f32(0.804801), f32(0.555656),
				f32(0.208671)],
			[f32(0.830847), f32(-0.06019), f32(-0.553237)],
			[f32(0.848333), f32(0.356899),
				f32(-0.391094)],
			[f32(0.946332), f32(-0.1508), f32(0.285859)],
			[f32(0.96289), f32(-0.22004), f32(-0.156284)],
			[f32(0.980377), f32(0.197049),
				f32(0.005858)]]
		faces:    [[30, 24, 37], [14, 28, 26], [11, 13, 22], [25, 38, 31],
			[48, 56, 55], [59, 57, 58], [39, 41, 50], [43, 49, 54],
			[40, 46, 34], [45, 36, 32], [53, 52, 44], [51, 42, 47],
			[21, 19, 10], [27, 15, 16], [33, 35, 23], [29, 20, 17],
			[18, 8, 12], [1, 3, 7], [5, 4, 0], [6, 9, 2], [18, 12, 24, 30],
			[24, 26, 39, 37], [26, 28, 41, 39], [11, 22, 28, 14],
			[13, 25, 31, 22], [31, 38, 49, 43], [30, 37, 48, 40],
			[56, 59, 58, 55], [58, 57, 52, 53], [50, 54, 59, 56],
			[41, 43, 54, 50], [49, 38, 42, 51], [48, 55, 46, 40],
			[46, 45, 32, 34], [36, 44, 33, 27], [53, 44, 36, 45],
			[57, 51, 47, 52], [47, 42, 29, 35], [34, 32, 19, 21],
			[19, 16, 5, 10], [16, 15, 4, 5], [33, 23, 15, 27],
			[35, 29, 17, 23], [17, 20, 9, 6], [21, 10, 8, 18],
			[8, 1, 7, 12], [7, 3, 11, 14], [0, 2, 3, 1], [4, 6, 2, 0],
			[9, 20, 25, 13], [12, 7, 14, 26, 24], [22, 31, 43, 41, 28],
			[37, 39, 50, 56, 48], [54, 49, 51, 57, 59], [55, 58, 53, 45, 46],
			[52, 47, 35, 33, 44], [32, 36, 27, 16, 19], [23, 17, 6, 4, 15],
			[10, 5, 0, 1, 8], [2, 9, 13, 11, 3], [18, 30, 40, 34, 21],
			[20, 29, 42, 38, 25]]
	},
	&Polyhedron{
		name:     'j76'
		vertexes: [[f32(-0.975594), f32(-0.152802), f32(-0.163647)],
			[f32(-0.930864), f32(0.290583), f32(-0.105382)],
			[f32(-0.885816), f32(-0.354103),
				f32(0.228021)],
			[f32(-0.840234), f32(-0.110417), f32(-0.590106)],
			[f32(-0.813441), f32(0.363309), f32(0.322296)],
			[f32(-0.812393), f32(-0.508854),
				f32(-0.384052)],
			[f32(-0.795504), f32(0.332968), f32(-0.531841)],
			[f32(-0.7856), f32(-0.035128),
				f32(0.52835)],
			[f32(-0.722614), f32(-0.710155), f32(0.007616)],
			[f32(-0.695288), f32(0.651943),
				f32(-0.231511)],
			[f32(-0.605191), f32(-0.637428), f32(0.435294)],
			[f32(-0.577865), f32(0.724669),
				f32(0.196167)],
			[f32(-0.531438), f32(-0.243136), f32(-0.888462)],
			[f32(-0.504975), f32(-0.318454), f32(0.735624)],
			[f32(-0.503596), f32(-0.641573),
				f32(-0.682408)],
			[f32(-0.488086), f32(0.523369), f32(0.587835)],
			[f32(-0.460245), f32(0.124931),
				f32(0.79389)],
			[f32(-0.459063), f32(0.474276), f32(-0.794187)],
			[f32(-0.358847), f32(0.793251),
				f32(-0.493857)],
			[f32(-0.358332), f32(-0.967284), f32(-0.048676)],
			[f32(-0.295861), f32(0.118224), f32(-1.01459)],
			[f32(-0.240909), f32(-0.894558),
				f32(0.379002)],
			[f32(-0.222972), f32(-0.924899), f32(-0.475135)],
			[f32(-0.168853), f32(0.910925), f32(0.19814)],
			[f32(-0.079074), f32(0.709624),
				f32(0.589809)],
			[f32(-0.078756), f32(-0.378446), f32(0.864946)],
			[f32(-0.050051), f32(0.660532),
				f32(-0.792214)],
			[f32(-0.034026), f32(0.064939), f32(0.923211)],
			[f32(-0.033492), f32(0.95331),
				f32(-0.228318)],
			[f32(0.067887), f32(-1.02728), f32(0.080646)],
			[f32(0.084446), f32(-0.734498),
				f32(0.644541)],
			[f32(0.113151), f32(0.30448), f32(-1.01262)],
			[f32(0.201551), f32(0.426299), f32(0.797082)],
			[f32(0.203247), f32(-0.984891),
				f32(-0.345813)],
			[f32(0.257366), f32(0.850932), f32(0.327462)],
			[f32(0.275304), f32(0.820591),
				f32(-0.526675)],
			[f32(0.330256), f32(-0.192191), f32(0.866919)],
			[f32(0.392727), f32(0.893318),
				f32(-0.098997)],
			[f32(0.393242), f32(-0.867217), f32(0.346185)],
			[f32(0.493458), f32(-0.548243),
				f32(0.646514)],
			[f32(0.537991), f32(0.567607), f32(0.534736)],
			[f32(0.53937), f32(0.244487),
				f32(-0.883296)],
			[f32(0.565833), f32(0.169169), f32(0.74079)],
			[f32(0.61226), f32(-0.798636), f32(-0.34384)],
			[f32(0.639586), f32(0.563462),
				f32(-0.582967)],
			[f32(0.729683), f32(-0.725909), f32(0.083838)],
			[f32(0.757009), f32(0.636188),
				f32(-0.155289)],
			[f32(0.819995), f32(-0.038838), f32(-0.676023)],
			[f32(0.829899), f32(-0.406935),
				f32(0.384168)],
			[f32(0.846787), f32(0.434888), f32(0.236379)],
			[f32(0.847836), f32(-0.437276),
				f32(-0.469969)],
			[f32(0.874629), f32(0.03645), f32(0.442434)],
			[f32(0.920211), f32(0.280136),
				f32(-0.375693)],
			[f32(0.965259), f32(-0.364549), f32(-0.042291)],
			[f32(1.00999), f32(0.078836),
				f32(0.015975)]]
		faces:    [[26, 17, 18], [6, 1, 9], [3, 5, 0], [8, 10, 2],
			[35, 28, 37], [23, 24, 34], [11, 4, 15], [7, 13, 16],
			[44, 46, 52], [49, 51, 54], [40, 32, 42], [27, 25, 36],
			[53, 48, 45], [39, 30, 38], [29, 21, 19], [31, 20, 17, 26],
			[17, 6, 9, 18], [9, 1, 4, 11], [3, 0, 1, 6], [5, 8, 2, 0],
			[2, 10, 13, 7], [26, 18, 28, 35], [28, 23, 34, 37],
			[34, 24, 32, 40], [11, 15, 24, 23], [4, 7, 16, 15],
			[16, 13, 25, 27], [35, 37, 46, 44], [46, 49, 54, 52],
			[54, 51, 48, 53], [40, 42, 51, 49], [32, 27, 36, 42],
			[36, 25, 30, 39], [44, 52, 47, 41], [53, 45, 43, 50],
			[48, 39, 38, 45], [38, 30, 21, 29], [12, 14, 5, 3],
			[33, 29, 19, 22], [19, 21, 10, 8], [20, 12, 3, 6, 17],
			[0, 2, 7, 4, 1], [18, 9, 11, 23, 28], [15, 16, 27, 32, 24],
			[37, 34, 40, 49, 46], [42, 36, 39, 48, 51], [52, 54, 53, 50, 47],
			[45, 38, 29, 33, 43], [22, 19, 8, 5, 14], [31, 26, 35, 44, 41],
			[21, 30, 25, 13, 10], [41, 47, 50, 43, 33, 22, 14, 12, 20, 31]]
	},
	&Polyhedron{
		name:     'j77'
		vertexes: [[f32(-0.965273), f32(-0.178368), f32(-0.195819)],
			[f32(-0.921193), f32(0.268836), f32(-0.202934)],
			[f32(-0.899923), f32(-0.317663),
				f32(0.226452)],
			[f32(-0.828599), f32(0.405929), f32(0.214939)],
			[f32(-0.815454), f32(0.043453),
				f32(0.480314)],
			[f32(-0.804857), f32(-0.20085), f32(-0.615041)],
			[f32(-0.791711), f32(-0.563327),
				f32(-0.349666)],
			[f32(-0.760776), f32(0.246354), f32(-0.622156)],
			[f32(-0.726361), f32(-0.702622),
				f32(0.072605)],
			[f32(-0.676307), f32(0.60747), f32(-0.368293)],
			[f32(-0.633767), f32(-0.565529),
				f32(0.490477)],
			[f32(-0.583713), f32(0.744563), f32(0.049579)],
			[f32(-0.582414), f32(0.411487),
				f32(0.590902)],
			[f32(-0.549298), f32(-0.204413), f32(0.74434)],
			[f32(-0.479947), f32(-0.376522),
				f32(-0.871086)],
			[f32(-0.466801), f32(-0.738998), f32(-0.605711)],
			[f32(-0.408623), f32(0.347071), f32(-0.882598)],
			[f32(-0.361062), f32(-0.964382),
				f32(0.077537)],
			[f32(-0.337528), f32(0.750121), f32(0.425542)],
			[f32(-0.324153), f32(0.708187),
				f32(-0.628736)],
			[f32(-0.316259), f32(0.163621), f32(0.854928)],
			[f32(-0.268468), f32(-0.827289),
				f32(0.49541)],
			[f32(-0.235061), f32(-0.037888), f32(-1.03645)],
			[f32(-0.200645), f32(-0.986864),
				f32(-0.341685)],
			[f32(-0.174334), f32(0.930008), f32(0.047397)],
			[f32(-0.131794), f32(-0.242991),
				f32(0.906168)],
			[f32(-0.013917), f32(0.907526), f32(-0.371825)],
			[f32(0.000756), f32(0.532515),
				f32(-0.88478)],
			[f32(0.041768), f32(-0.62795), f32(0.752321)],
			[f32(0.056442), f32(-1.00296),
				f32(0.239365)],
			[f32(0.079975), f32(0.711542), f32(0.58737)],
			[f32(0.093121), f32(0.349066), f32(0.852745)],
			[f32(0.174319), f32(0.147557),
				f32(-1.03863)],
			[f32(0.216858), f32(-1.02544), f32(-0.179857)],
			[f32(0.24317), f32(0.89143), f32(0.209225)],
			[f32(0.277585), f32(-0.057546), f32(0.903985)],
			[f32(0.310993), f32(0.731855),
				f32(-0.62787)],
			[f32(0.366678), f32(-0.803621), f32(0.496276)],
			[f32(0.403586), f32(0.868948),
				f32(-0.209997)],
			[f32(0.451147), f32(-0.442505), f32(0.750138)],
			[f32(0.509326), f32(0.643564),
				f32(0.473251)],
			[f32(0.522471), f32(0.281088), f32(0.738626)],
			[f32(0.591822), f32(0.108979), f32(-0.8768)],
			[f32(0.626237), f32(-0.839998),
				f32(-0.182039)],
			[f32(0.676292), f32(0.470095), f32(-0.622937)],
			[f32(0.718831), f32(-0.702904),
				f32(0.235834)],
			[f32(0.768885), f32(0.607188), f32(-0.205064)],
			[f32(0.8033), f32(-0.341788),
				f32(0.489696)],
			[f32(0.834235), f32(0.467893), f32(0.217206)],
			[f32(0.847381), f32(0.105416),
				f32(0.482581)],
			[f32(0.857978), f32(-0.138887), f32(-0.612774)],
			[f32(0.871123), f32(-0.501364),
				f32(-0.347399)],
			[f32(0.942447), f32(0.222229), f32(-0.358911)],
			[f32(0.963717), f32(-0.36427),
				f32(0.070474)],
			[f32(1.0078), f32(0.082934), f32(0.063359)]]
		faces:    [[27, 16, 19], [7, 1, 9], [5, 6, 0], [8, 10, 2],
			[36, 26, 38], [11, 18, 24], [3, 4, 12], [13, 25, 20],
			[44, 46, 52], [48, 49, 54], [34, 30, 40], [31, 35, 41],
			[53, 47, 45], [39, 28, 37], [29, 21, 17], [32, 22, 16, 27],
			[16, 7, 9, 19], [9, 1, 3, 11], [5, 0, 1, 7], [6, 8, 2, 0],
			[2, 10, 13, 4], [27, 19, 26, 36], [26, 24, 34, 38],
			[24, 18, 30, 34], [3, 12, 18, 11], [4, 13, 20, 12],
			[20, 25, 35, 31], [36, 38, 46, 44], [46, 48, 54, 52],
			[54, 49, 47, 53], [40, 41, 49, 48], [30, 31, 41, 40],
			[35, 25, 28, 39], [44, 52, 50, 42], [53, 45, 43, 51],
			[47, 39, 37, 45], [37, 28, 21, 29], [14, 15, 6, 5],
			[33, 29, 17, 23], [17, 21, 10, 8], [22, 14, 5, 7, 16],
			[0, 2, 4, 3, 1], [19, 9, 11, 24, 26], [12, 20, 31, 30, 18],
			[38, 34, 40, 48, 46], [41, 35, 39, 47, 49], [52, 54, 53, 51, 50],
			[45, 37, 29, 33, 43], [23, 17, 8, 6, 15], [32, 27, 36, 44, 42],
			[21, 28, 25, 13, 10], [42, 50, 51, 43, 33, 23, 15, 14, 22, 32]]
	},
	&Polyhedron{
		name:     'j78'
		vertexes: [[f32(-0.969175), f32(0.215371), f32(-0.127391)],
			[f32(-0.952173), f32(-0.166819), f32(-0.363246)],
			[f32(-0.946899), f32(-0.019645), f32(0.255045)],
			[f32(-0.929897), f32(-0.401835),
				f32(0.01919)],
			[f32(-0.840084), f32(0.222491), f32(-0.557822)],
			[f32(-0.781766), f32(-0.392789),
				f32(0.443408)],
			[f32(-0.765536), f32(0.610272), f32(-0.059785)],
			[f32(-0.729493), f32(0.230008),
				f32(0.559009)],
			[f32(-0.721025), f32(-0.390315), f32(-0.677262)],
			[f32(-0.684982), f32(-0.770578), f32(-0.058468)],
			[f32(-0.636445), f32(0.617392), f32(-0.490216)],
			[f32(-0.617404), f32(0.619318),
				f32(0.364433)],
			[f32(-0.608936), f32(-0.001005), f32(-0.871838)],
			[f32(-0.56436), f32(-0.143136), f32(0.747372)],
			[f32(-0.555892), f32(-0.763458),
				f32(-0.488899)],
			[f32(-0.536851), f32(-0.761533), f32(0.36575)],
			[f32(-0.419039), f32(0.867044),
				f32(-0.186253)],
			[f32(-0.360721), f32(0.251764), f32(0.814977)],
			[f32(-0.305703), f32(-0.985028),
				f32(0.051734)],
			[f32(-0.279442), f32(0.637958), f32(-0.76245)],
			[f32(-0.270908), f32(0.87609),
				f32(0.237966)],
			[f32(-0.26244), f32(0.255768), f32(-0.998305)],
			[f32(-0.248632), f32(0.641074),
				f32(0.620402)],
			[f32(-0.185081), f32(-0.357586), f32(0.857574)],
			[f32(-0.176613), f32(-0.977908),
				f32(-0.378698)],
			[f32(-0.168079), f32(-0.739776), f32(0.621718)],
			[f32(-0.062036), f32(0.887611),
				f32(-0.458486)],
			[f32(0.018558), f32(0.037315), f32(0.925179)],
			[f32(0.063069), f32(-0.963271),
				f32(0.307702)],
			[f32(0.169112), f32(0.664116), f32(-0.772503)],
			[f32(0.177646), f32(0.902248),
				f32(0.227913)],
			[f32(0.186114), f32(0.281925), f32(-1.00836)],
			[f32(0.199922), f32(0.667232),
				f32(0.610349)],
			[f32(0.211888), f32(-0.546211), f32(0.763647)],
			[f32(0.271941), f32(-0.951751),
				f32(-0.38875)],
			[f32(0.306736), f32(0.909368), f32(-0.202518)],
			[f32(0.365054), f32(0.294088),
				f32(0.798712)],
			[f32(0.415527), f32(-0.151311), f32(0.831252)],
			[f32(0.420072), f32(-0.942705),
				f32(0.035468)],
			[f32(0.443036), f32(-0.769707), f32(0.44963)],
			[f32(0.537884), f32(0.685872),
				f32(-0.516534)],
			[f32(0.556925), f32(0.687798), f32(0.338115)],
			[f32(0.565393), f32(0.067476),
				f32(-0.898156)],
			[f32(0.618437), f32(-0.694978), f32(-0.515217)],
			[f32(0.686015), f32(0.694918),
				f32(-0.092316)],
			[f32(0.722058), f32(0.314654), f32(0.526478)],
			[f32(0.730526), f32(-0.305668),
				f32(-0.709793)],
			[f32(0.766569), f32(-0.685932), f32(-0.090999)],
			[f32(0.77253), f32(-0.130744),
				f32(0.559019)],
			[f32(0.782799), f32(0.317129), f32(-0.594192)],
			[f32(0.789532), f32(-0.512934),
				f32(0.323163)],
			[f32(0.93093), f32(0.326175), f32(-0.169974)],
			[f32(0.947932), f32(-0.056015),
				f32(-0.405829)],
			[f32(0.953206), f32(0.091159), f32(0.212462)],
			[f32(0.970208), f32(-0.291031),
				f32(-0.023393)]]
		faces:    [[29, 19, 26], [10, 6, 16], [4, 1, 0], [3, 5, 2],
			[40, 35, 44], [30, 32, 41], [20, 11, 22], [7, 13, 17],
			[49, 51, 52], [45, 48, 53], [36, 27, 37], [23, 25, 33],
			[54, 50, 47], [39, 28, 38], [18, 15, 9], [31, 21, 19, 29],
			[19, 10, 16, 26], [16, 6, 11, 20], [4, 0, 6, 10],
			[1, 3, 2, 0], [2, 5, 13, 7], [29, 26, 35, 40], [35, 30, 41, 44],
			[41, 32, 36, 45], [20, 22, 32, 30], [11, 7, 17, 22],
			[17, 13, 23, 27], [40, 44, 51, 49], [51, 53, 54, 52],
			[53, 48, 50, 54], [36, 37, 48, 45], [27, 23, 33, 37],
			[33, 25, 28, 39], [49, 52, 46, 42], [47, 38, 34, 43],
			[50, 39, 38, 47], [28, 25, 15, 18], [12, 8, 1, 4],
			[24, 18, 9, 14], [9, 15, 5, 3], [21, 12, 4, 10, 19],
			[0, 2, 7, 11, 6], [26, 16, 20, 30, 35], [22, 17, 27, 36, 32],
			[44, 41, 45, 53, 51], [37, 33, 39, 50, 48], [52, 54, 47, 43, 46],
			[38, 28, 18, 24, 34], [14, 9, 3, 1, 8], [31, 29, 40, 49, 42],
			[15, 25, 23, 13, 5], [42, 46, 43, 34, 24, 14, 8, 12, 21, 31]]
	},
	&Polyhedron{
		name:     'j79'
		vertexes: [[f32(-1.03566), f32(0.17951), f32(0.161516)],
			[f32(-1.02789), f32(0.048482), f32(-0.268318)],
			[f32(-0.891113), f32(0.078842),
				f32(0.574986)],
			[f32(-0.870771), f32(-0.264193), f32(-0.550334)],
			[f32(-0.833419), f32(0.579967), f32(0.188311)],
			[f32(-0.820848), f32(0.367959),
				f32(-0.507174)],
			[f32(-0.700657), f32(0.696435), f32(-0.224962)],
			[f32(-0.68887), f32(0.479299),
				f32(0.601781)],
			[f32(-0.663727), f32(0.055284), f32(-0.78919)],
			[f32(-0.649458), f32(-0.215069),
				f32(0.814161)],
			[f32(-0.624314), f32(-0.639084), f32(-0.576811)],
			[f32(-0.485083), f32(0.858791), f32(0.134418)],
			[f32(-0.461483), f32(0.455741),
				f32(-0.762395)],
			[f32(-0.403), f32(-0.58996), f32(0.787683)],
			[f32(-0.382659), f32(-0.932996),
				f32(-0.337637)],
			[f32(-0.341293), f32(0.784217), f32(-0.480183)],
			[f32(-0.340534), f32(0.758124),
				f32(0.547888)],
			[f32(-0.322222), f32(0.432884), f32(0.857516)],
			[f32(-0.297863), f32(0.00374),
				f32(0.988774)],
			[f32(-0.289308), f32(-0.122159), f32(-0.96329)],
			[f32(-0.26495), f32(-0.551303),
				f32(-0.832032)],
			[f32(-0.245879), f32(-0.902636), f32(0.505667)],
			[f32(-0.238109), f32(-1.03366),
				f32(0.075833)],
			[f32(-0.125719), f32(0.946573), f32(-0.120803)],
			[f32(-0.087065), f32(0.278298),
				f32(-0.936494)],
			[f32(-0.051406), f32(-0.371151), f32(0.962296)],
			[f32(-0.023294), f32(-0.845214),
				f32(-0.592857)],
			[f32(0.107408), f32(0.809782), f32(-0.479865)],
			[f32(0.108167), f32(0.783689),
				f32(0.548206)],
			[f32(0.110226), f32(-0.32589), f32(-0.934099)],
			[f32(0.126479), f32(0.458449),
				f32(0.857834)],
			[f32(0.150837), f32(0.029306), f32(0.989092)],
			[f32(0.202822), f32(-0.87707),
				f32(0.505985)],
			[f32(0.210592), f32(-1.0081), f32(0.076151)],
			[f32(0.24093), f32(0.900157), f32(0.134932)],
			[f32(0.264529), f32(0.497107),
				f32(-0.761881)],
			[f32(0.312469), f32(0.074567), f32(-0.907304)],
			[f32(0.323013), f32(-0.548594),
				f32(0.788197)],
			[f32(0.343354), f32(-0.89163), f32(-0.337123)],
			[f32(0.351882), f32(-0.619801),
				f32(-0.694925)],
			[f32(0.474057), f32(0.763367), f32(-0.224131)],
			[f32(0.485843), f32(0.546231),
				f32(0.602613)],
			[f32(0.525256), f32(-0.148138), f32(0.814992)],
			[f32(0.562186), f32(-0.789288),
				f32(0.250764)],
			[f32(0.618606), f32(0.662699), f32(0.189339)],
			[f32(0.631178), f32(0.450691),
				f32(-0.506147)],
			[f32(0.679118), f32(0.028151), f32(-0.651569)],
			[f32(0.682377), f32(-0.460813),
				f32(0.532976)],
			[f32(0.694949), f32(-0.672821), f32(-0.16251)],
			[f32(0.703476), f32(-0.400992),
				f32(-0.520312)],
			[f32(0.7323), f32(0.17134), f32(0.576135)], [f32(0.865063), f32(0.287808), f32(0.162862)],
			[f32(0.872833), f32(0.15678), f32(-0.266972)],
			[f32(0.889422), f32(-0.141336),
				f32(0.29412)],
			[f32(0.897192), f32(-0.272364), f32(-0.135714)]]
		faces:    [[7, 17, 16], [30, 41, 28], [18, 25, 31], [37, 47, 42],
			[4, 11, 6], [23, 27, 15], [34, 44, 40], [50, 53, 51],
			[5, 12, 8], [35, 36, 24], [45, 52, 46], [54, 48, 49],
			[19, 29, 20], [39, 38, 26], [33, 43, 32], [0, 2, 7, 4],
			[17, 30, 28, 16], [28, 41, 44, 34], [18, 31, 30, 17],
			[25, 37, 42, 31], [42, 47, 53, 50], [7, 16, 11, 4],
			[11, 23, 15, 6], [27, 40, 45, 35], [34, 40, 27, 23],
			[41, 50, 51, 44], [51, 53, 54, 52], [6, 15, 12, 5],
			[12, 24, 19, 8], [24, 36, 29, 19], [45, 46, 36, 35],
			[52, 54, 49, 46], [49, 48, 38, 39], [5, 8, 3, 1],
			[20, 26, 14, 10], [29, 39, 26, 20], [38, 48, 43, 33],
			[9, 13, 25, 18], [22, 33, 32, 21], [32, 43, 47, 37],
			[2, 9, 18, 17, 7], [31, 42, 50, 41, 30], [16, 28, 34, 23, 11],
			[44, 51, 52, 45, 40], [15, 27, 35, 24, 12], [46, 49, 39, 29, 36],
			[8, 19, 20, 10, 3], [26, 38, 33, 22, 14], [21, 32, 37, 25, 13],
			[0, 4, 6, 5, 1], [43, 48, 54, 53, 47], [1, 3, 10, 14, 22, 21, 13, 9, 2, 0]]
	},
	&Polyhedron{
		name:     'j80'
		vertexes: [[f32(-0.981435), f32(-0.157408), f32(-0.109585)],
			[f32(-0.942153), f32(-0.069788), f32(0.327838)],
			[f32(-0.91551), f32(0.22466),
				f32(-0.333721)],
			[f32(-0.85195), f32(0.366431), f32(0.374044)],
			[f32(-0.835484), f32(0.54841),
				f32(-0.034822)],
			[f32(-0.80426), f32(-0.38784), f32(-0.450273)],
			[f32(-0.738335), f32(-0.005772),
				f32(-0.67441)],
			[f32(-0.701418), f32(-0.15845), f32(0.694914)],
			[f32(-0.648132), f32(0.430447),
				f32(-0.628204)],
			[f32(-0.611216), f32(0.27777), f32(0.74112)],
			[f32(-0.568107), f32(0.754197),
				f32(-0.329305)],
			[f32(-0.545291), f32(0.659837), f32(0.516984)],
			[f32(-0.528825), f32(0.841816),
				f32(0.108118)],
			[f32(-0.478303), f32(-0.673069), f32(-0.564096)],
			[f32(-0.371634), f32(-0.05487), f32(-0.926756)],
			[f32(-0.351184), f32(-0.389527),
				f32(0.851433)],
			[f32(-0.281432), f32(0.381349), f32(-0.88055)],
			[f32(-0.210926), f32(-0.467282),
				f32(-0.858579)],
			[f32(-0.205234), f32(0.316291), f32(0.926196)],
			[f32(-0.151948), f32(0.905188),
				f32(-0.396922)],
			[f32(-0.139309), f32(0.698359), f32(0.70206)],
			[f32(-0.128068), f32(-0.904145),
				f32(-0.407577)],
			[f32(-0.112666), f32(0.992807), f32(0.040501)],
			[f32(-0.044525), f32(-0.09612),
				f32(0.994373)],
			[f32(-0.025227), f32(-0.674755), f32(0.73761)],
			[f32(0.025227), f32(0.674755),
				f32(-0.73761)],
			[f32(0.044525), f32(0.096121), f32(-0.994373)],
			[f32(0.112666), f32(-0.992807),
				f32(-0.040501)],
			[f32(0.128068), f32(0.904146), f32(0.407577)],
			[f32(0.139309), f32(-0.698358),
				f32(-0.70206)],
			[f32(0.151948), f32(-0.905188), f32(0.396922)],
			[f32(0.205234), f32(-0.316291),
				f32(-0.926196)],
			[f32(0.210926), f32(0.467282), f32(0.858579)],
			[f32(0.281432), f32(-0.381349),
				f32(0.88055)],
			[f32(0.351184), f32(0.389527), f32(-0.851433)],
			[f32(0.371634), f32(0.05487),
				f32(0.926756)],
			[f32(0.478303), f32(0.673069), f32(0.564096)],
			[f32(0.528825), f32(-0.841816),
				f32(-0.108118)],
			[f32(0.545291), f32(-0.659837), f32(-0.516984)],
			[f32(0.568107), f32(-0.754197),
				f32(0.329305)],
			[f32(0.611216), f32(-0.277769), f32(-0.74112)],
			[f32(0.648133), f32(-0.430447),
				f32(0.628204)],
			[f32(0.701419), f32(0.15845), f32(-0.694914)],
			[f32(0.738335), f32(0.005773), f32(0.67441)],
			[f32(0.80426), f32(0.387841), f32(0.450273)],
			[f32(0.835484), f32(-0.54841), f32(0.034822)],
			[f32(0.85195), f32(-0.366431),
				f32(-0.374044)],
			[f32(0.91551), f32(-0.22466), f32(0.333721)],
			[f32(0.942153), f32(0.069789),
				f32(-0.327838)],
			[f32(0.981435), f32(0.157408), f32(0.109585)]]
		faces:    [[12, 10, 4], [8, 6, 2], [16, 26, 14], [31, 29, 17],
			[11, 3, 9], [20, 18, 32], [23, 33, 35], [43, 41, 47],
			[39, 37, 45], [46, 38, 40], [22, 19, 10, 12], [10, 8, 2, 4],
			[2, 6, 5, 0], [16, 14, 6, 8], [26, 31, 17, 14], [17, 29, 21, 13],
			[12, 4, 3, 11], [3, 1, 7, 9], [11, 9, 18, 20], [18, 23, 35, 32],
			[35, 33, 41, 43], [15, 24, 33, 23], [30, 27, 37, 39],
			[20, 32, 36, 28], [43, 47, 49, 44], [41, 39, 45, 47],
			[45, 37, 38, 46], [25, 34, 26, 16], [48, 46, 40, 42],
			[40, 38, 29, 31], [19, 25, 16, 8, 10], [14, 17, 13, 5, 6],
			[4, 2, 0, 1, 3], [9, 7, 15, 23, 18], [24, 30, 39, 41, 33],
			[32, 35, 43, 44, 36], [47, 45, 46, 48, 49], [42, 40, 31, 26, 34],
			[22, 12, 11, 20, 28], [38, 37, 27, 21, 29], [24, 15, 7, 1, 0, 5, 13, 21, 27, 30],
			[28, 36, 44, 49, 48, 42, 34, 25, 19, 22]]
	},
	&Polyhedron{
		name:     'j81'
		vertexes: [[f32(-0.91554), f32(-0.17156), f32(0.190699)],
			[f32(-0.874123), f32(-0.21861), f32(-0.254883)],
			[f32(-0.873513), f32(0.274357),
				f32(0.14752)],
			[f32(-0.832096), f32(0.227307), f32(-0.298062)],
			[f32(-0.790984), f32(-0.567471),
				f32(0.016881)],
			[f32(-0.738991), f32(-0.290113), f32(0.587244)],
			[f32(-0.680957), f32(0.599954),
				f32(-0.096163)],
			[f32(-0.670991), f32(0.431396), f32(0.517379)],
			[f32(-0.630562), f32(-0.413291),
				f32(-0.579305)],
			[f32(-0.614436), f32(-0.686024), f32(0.413427)],
			[f32(-0.587852), f32(0.082534),
				f32(0.789144)],
			[f32(-0.562561), f32(0.308217), f32(-0.64917)],
			[f32(-0.547423), f32(-0.762153),
				f32(-0.30754)],
			[f32(-0.478435), f32(0.756993), f32(0.273697)],
			[f32(-0.438006), f32(-0.087694),
				f32(-0.822987)],
			[f32(-0.411421), f32(0.680864), f32(-0.44727)],
			[f32(-0.301886), f32(0.63844),
				f32(0.670242)],
			[f32(-0.277887), f32(-0.681242), f32(-0.658648)],
			[f32(-0.261761), f32(-0.953976), f32(0.334084)],
			[f32(-0.220345), f32(-1.00103),
				f32(-0.111498)],
			[f32(-0.218747), f32(0.289578), f32(0.942007)],
			[f32(-0.16786), f32(0.486183),
				f32(-0.771692)],
			[f32(-0.085331), f32(-0.355646), f32(-0.90233)],
			[f32(-0.083733), f32(0.934958),
				f32(0.151175)],
			[f32(-0.043304), f32(0.090271), f32(-0.945509)],
			[f32(-0.042317), f32(0.887908),
				f32(-0.294407)],
			[f32(0.049191), f32(-0.920115), f32(-0.462606)],
			[f32(0.092815), f32(0.816405),
				f32(0.54772)],
			[f32(0.184323), f32(-0.991618), f32(0.379522)],
			[f32(0.201245), f32(0.693227),
				f32(-0.618829)],
			[f32(0.225739), f32(-1.03867), f32(-0.06606)],
			[f32(0.227337), f32(0.251936),
				f32(0.987445)],
			[f32(0.360753), f32(-0.393288), f32(-0.856892)],
			[f32(0.362351), f32(0.897316),
				f32(0.196613)],
			[f32(0.40278), f32(0.052629), f32(-0.900071)],
			[f32(0.403767), f32(0.850266),
				f32(-0.24897)],
			[f32(0.419893), f32(0.577533), f32(0.743762)],
			[f32(0.443892), f32(-0.74215),
				f32(-0.585128)],
			[f32(0.553427), f32(-0.784574), f32(0.532385)],
			[f32(0.553919), f32(0.425276),
				f32(-0.698172)],
			[f32(0.580011), f32(-0.016016), f32(0.908102)],
			[f32(0.62044), f32(-0.860702),
				f32(-0.188582)],
			[f32(0.689428), f32(0.658443), f32(0.392655)],
			[f32(0.704567), f32(-0.411927),
				f32(0.734284)],
			[f32(0.756442), f32(0.582315), f32(-0.328312)],
			[f32(0.772567), f32(0.309582),
				f32(0.664419)],
			[f32(0.822963), f32(-0.703664), f32(0.181277)],
			[f32(0.93299), f32(0.463762),
				f32(0.068233)],
			[f32(0.974102), f32(-0.331017), f32(0.383177)],
			[f32(1.01613), f32(0.1149), f32(0.339998)]]
		faces:    [[35, 29, 25], [21, 11, 15], [24, 22, 14], [17, 12, 8],
			[33, 23, 27], [13, 7, 16], [6, 3, 2], [1, 4, 0], [42, 36, 45],
			[30, 19, 26], [44, 39, 29, 35], [29, 21, 15, 25],
			[15, 11, 3, 6], [24, 14, 11, 21], [22, 17, 8, 14],
			[8, 12, 4, 1], [35, 25, 23, 33], [23, 13, 16, 27],
			[16, 7, 10, 20], [6, 2, 7, 13], [3, 1, 0, 2], [0, 4, 9, 5],
			[33, 27, 36, 42], [36, 31, 40, 45], [42, 45, 49, 47],
			[43, 38, 46, 48], [28, 18, 19, 30], [34, 32, 22, 24],
			[41, 30, 26, 37], [26, 19, 12, 17], [39, 34, 24, 21, 29],
			[14, 8, 1, 3, 11], [25, 15, 6, 13, 23], [2, 0, 5, 10, 7],
			[27, 16, 20, 31, 36], [45, 40, 43, 48, 49], [38, 28, 30, 41, 46],
			[37, 26, 17, 22, 32], [44, 35, 33, 42, 47], [19, 18, 9, 4, 12],
			[38, 43, 40, 31, 20, 10, 5, 9, 18, 28], [47, 49, 48, 46, 41, 37, 32, 34, 39, 44]]
	},
	&Polyhedron{
		name:     'j82'
		vertexes: [[f32(-0.915244), f32(-0.149547), f32(0.004878)],
			[f32(-0.857812), f32(0.261033), f32(-0.170045)],
			[f32(-0.853796), f32(0.017864),
				f32(0.418001)],
			[f32(-0.796364), f32(0.428444), f32(0.243078)],
			[f32(-0.772518), f32(-0.333547),
				f32(-0.380149)],
			[f32(-0.759676), f32(-0.571754), f32(0.001381)],
			[f32(-0.715086), f32(0.077033),
				f32(-0.555071)],
			[f32(-0.660252), f32(-0.300878), f32(0.669827)],
			[f32(-0.638771), f32(0.334916),
				f32(0.65404)],
			[f32(-0.609317), f32(0.503159), f32(-0.456572)],
			[f32(-0.602083), f32(-0.665282),
				f32(0.412342)],
			[f32(-0.509893), f32(0.774035), f32(0.211875)],
			[f32(-0.463372), f32(-0.606112),
				f32(-0.56073)],
			[f32(-0.45053), f32(-0.844319), f32(-0.1792)],
			[f32(-0.445227), f32(0.016174),
				f32(0.905866)],
			[f32(-0.394292), f32(0.820211), f32(-0.220533)],
			[f32(-0.370445), f32(0.05822),
				f32(-0.84376)],
			[f32(-0.3523), f32(0.680507), f32(0.622836)],
			[f32(-0.292937), f32(-0.937847),
				f32(0.231761)],
			[f32(-0.264676), f32(0.484346), f32(-0.745261)],
			[f32(-0.214877), f32(-0.363987),
				f32(-0.847257)],
			[f32(-0.105889), f32(-0.863132), f32(-0.467889)],
			[f32(-0.103806), f32(0.922633), f32(0.336308)],
			[f32(-0.049651), f32(0.801399),
				f32(-0.509222)],
			[f32(-0.039139), f32(0.164772), f32(1.0303)],
			[f32(0.011796), f32(0.968809),
				f32(-0.096099)],
			[f32(0.018293), f32(0.575352), f32(0.855378)],
			[f32(0.04447), f32(0.211781),
				f32(-0.925842)],
			[f32(0.142605), f32(-0.621006), f32(-0.754417)],
			[f32(0.149102), f32(-1.01446),
				f32(0.197061)],
			[f32(0.200037), f32(-0.210426), f32(-0.929339)],
			[f32(0.264704), f32(-0.968287),
				f32(-0.235347)],
			[f32(0.266787), f32(0.817478), f32(0.56885)],
			[f32(0.392388), f32(0.724782),
				f32(-0.543923)],
			[f32(0.4029), f32(0.088156), f32(0.9956)], [f32(0.450558), f32(0.360379), f32(-0.801408)],
			[f32(0.453835), f32(0.892193), f32(-0.1308)],
			[f32(0.460331), f32(0.498736), f32(0.820677)],
			[f32(0.513198), f32(-0.726161),
				f32(-0.521875)],
			[f32(0.55519), f32(-0.865866), f32(0.321494)],
			[f32(0.606125), f32(-0.061828),
				f32(-0.804905)],
			[f32(0.611428), f32(0.798665), f32(0.280161)],
			[f32(0.670792), f32(-0.819689),
				f32(-0.110913)],
			[f32(0.712045), f32(-0.18441), f32(0.815019)],
			[f32(0.770215), f32(-0.548813),
				f32(0.557534)],
			[f32(0.799669), f32(-0.38057), f32(-0.553078)],
			[f32(0.804972), f32(0.479923),
				f32(0.531988)],
			[f32(0.957263), f32(-0.474098), f32(-0.142117)],
			[f32(0.96054), f32(0.057716),
				f32(0.528491)],
			[f32(1.01871), f32(-0.306688), f32(0.271006)]]
		faces:    [[25, 23, 15], [27, 16, 19], [30, 28, 20], [21, 13, 12],
			[22, 11, 17], [3, 2, 8], [9, 6, 1], [4, 5, 0], [32, 26, 37],
			[42, 31, 38], [36, 33, 23, 25], [23, 19, 9, 15], [19, 16, 6, 9],
			[30, 20, 16, 27], [28, 21, 12, 20], [12, 13, 5, 4],
			[25, 15, 11, 22], [11, 3, 8, 17], [8, 2, 7, 14], [1, 0, 2, 3],
			[6, 4, 0, 1], [5, 13, 18, 10], [22, 17, 26, 32], [26, 24, 34, 37],
			[32, 37, 46, 41], [43, 44, 49, 48], [39, 29, 31, 42],
			[35, 40, 30, 27], [47, 42, 38, 45], [38, 31, 21, 28],
			[33, 35, 27, 19, 23], [20, 12, 4, 6, 16], [15, 9, 1, 3, 11],
			[0, 5, 10, 7, 2], [17, 8, 14, 24, 26], [37, 34, 43, 48, 46],
			[44, 39, 42, 47, 49], [45, 38, 28, 30, 40], [36, 25, 22, 32, 41],
			[31, 29, 18, 13, 21], [44, 43, 34, 24, 14, 7, 10, 18, 29, 39],
			[41, 46, 48, 49, 47, 45, 40, 35, 33, 36]]
	},
	&Polyhedron{
		name:     'j83'
		vertexes: [[f32(-0.932936), f32(0.189273), f32(0.192295)],
			[f32(-0.922398), f32(0.241407), f32(-0.253129)],
			[f32(-0.911995), f32(-0.249962),
				f32(0.280987)],
			[f32(-0.894943), f32(-0.165606), f32(-0.439724)],
			[f32(-0.888514), f32(-0.469289), f32(-0.109623)],
			[f32(-0.719187), f32(0.580372), f32(0.243128)],
			[f32(-0.712758), f32(0.27669),
				f32(0.57323)],
			[f32(-0.708649), f32(0.632507), f32(-0.202295)],
			[f32(-0.691817), f32(-0.162545),
				f32(0.661922)],
			[f32(-0.636773), f32(-0.433068), f32(-0.690809)],
			[f32(-0.630343), f32(-0.736751), f32(-0.360707)],
			[f32(-0.352393), f32(0.77395), f32(0.41407)],
			[f32(-0.345964), f32(0.470268),
				f32(0.744172)],
			[f32(-0.335341), f32(0.858306), f32(-0.306641)],
			[f32(-0.31208), f32(-0.240428),
				f32(0.887678)],
			[f32(-0.246498), f32(-0.458817), f32(-0.910477)],
			[f32(-0.236095), f32(-0.950186), f32(-0.376361)],
			[f32(-0.115163), f32(0.945723), f32(0.074294)],
			[f32(-0.098331), f32(0.150671),
				f32(0.938511)],
			[f32(0.001135), f32(-0.778414), f32(-0.716137)],
			[f32(0.027344), f32(0.696067),
				f32(0.639826)],
			[f32(0.054934), f32(0.832556), f32(-0.526309)],
			[f32(0.082168), f32(-0.453864),
				f32(0.872024)],
			[f32(0.12681), f32(-0.233018), f32(-1.01482)],
			[f32(0.143641), f32(-1.02807),
				f32(-0.150605)],
			[f32(0.264573), f32(0.867839), f32(0.30005)],
			[f32(0.274976), f32(0.37647), f32(0.834165)],
			[f32(0.275112), f32(0.919973),
				f32(-0.145374)],
			[f32(0.295917), f32(-0.062764), f32(0.922857)],
			[f32(0.313104), f32(0.565095),
				f32(-0.777393)],
			[f32(0.340339), f32(-0.721326), f32(0.620939)],
			[f32(0.340559), f32(0.158081),
				f32(-0.963989)],
			[f32(0.36382), f32(-0.940653), f32(0.23033)],
			[f32(0.374442), f32(-0.552615),
				f32(-0.820483)],
			[f32(0.380871), f32(-0.856297), f32(-0.490381)],
			[f32(0.658822), f32(0.654404),
				f32(0.284396)],
			[f32(0.665251), f32(0.350721), f32(0.614498)],
			[f32(0.66936), f32(0.706538),
				f32(-0.161028)],
			[f32(0.686192), f32(-0.088513), f32(0.703189)],
			[f32(0.692841), f32(0.487211),
				f32(-0.551637)],
			[f32(0.713646), f32(-0.495527), f32(0.516594)],
			[f32(0.720295), f32(0.080198),
				f32(-0.738233)],
			[f32(0.737127), f32(-0.714854), f32(0.125984)],
			[f32(0.741236), f32(-0.359037),
				f32(-0.649541)],
			[f32(0.747665), f32(-0.662719), f32(-0.31944)]]
		faces:    [[25, 27, 17], [20, 11, 12], [5, 0, 6], [26, 18, 28],
			[34, 19, 33], [35, 37, 27, 25], [27, 21, 13, 17],
			[25, 17, 11, 20], [11, 5, 6, 12], [6, 0, 2, 8], [7, 1, 0, 5],
			[3, 9, 10, 4], [20, 12, 18, 26], [18, 14, 22, 28],
			[26, 28, 38, 36], [30, 32, 42, 40], [24, 16, 19, 34],
			[39, 41, 31, 29], [44, 34, 33, 43], [33, 19, 15, 23],
			[37, 39, 29, 21, 27], [17, 13, 7, 5, 11], [1, 3, 4, 2, 0],
			[12, 6, 8, 14, 18], [28, 22, 30, 40, 38], [32, 24, 34, 44, 42],
			[43, 33, 23, 31, 41], [35, 25, 20, 26, 36], [19, 16, 10, 9, 15],
			[1, 7, 13, 21, 29, 31, 23, 15, 9, 3], [32, 30, 22, 14, 8, 2, 4, 10, 16, 24],
			[36, 38, 40, 42, 44, 43, 41, 39, 37, 35]]
	},
	&Polyhedron{
		name:     'j84'
		vertexes: [[f32(-0.768016), f32(0.559678), f32(0.635844)],
			[f32(-0.720709), f32(-0.093633), f32(-0.405339)],
			[f32(-0.6358), f32(-0.662351), f32(0.681929)],
			[f32(0.09848), f32(0.800885),
				f32(-0.202562)],
			[f32(0.269587), f32(-0.77416), f32(-0.143135)],
			[f32(0.285934), f32(-0.010665),
				f32(-1.1073)],
			[f32(0.352377), f32(0.066396), f32(0.750712)],
			[f32(1.11815), f32(0.11385), f32(-0.210152)]]
		faces:    [[6, 7, 3], [3, 7, 5], [3, 5, 1], [4, 7, 6],
			[7, 4, 5], [5, 4, 1], [4, 2, 1], [1, 2, 0], [1, 0, 3],
			[6, 2, 4], [2, 6, 0], [0, 6, 3]]
	},
	&Polyhedron{
		name:     'j85'
		vertexes: [[f32(-0.984789), f32(0.388776), f32(-0.318546)],
			[f32(-0.905986), f32(-0.50645), f32(-0.380955)],
			[f32(-0.774402), f32(-0.096785),
				f32(0.410496)],
			[f32(-0.648503), f32(0.795226), f32(0.411689)],
			[f32(-0.32762), f32(0.028199),
				f32(-0.818195)],
			[f32(-0.278924), f32(-0.81528), f32(0.187334)],
			[f32(-0.177548), f32(0.78687),
				f32(-0.356208)],
			[f32(-0.134682), f32(-0.843968), f32(-0.701432)],
			[f32(-0.06669), f32(0.257644), f32(0.840681)],
			[f32(0.229454), f32(0.996879),
				f32(0.419536)],
			[f32(0.428788), f32(-0.460851), f32(0.617519)],
			[f32(0.523163), f32(-0.229235),
				f32(-0.671807)],
			[f32(0.55373), f32(-0.948137), f32(-0.129793)],
			[f32(0.673235), f32(0.529435),
				f32(-0.20982)],
			[f32(0.811213), f32(0.353538), f32(0.662851)],
			[f32(1.07956), f32(-0.235865), f32(0.03665)]]
		faces:    [[13, 9, 14], [9, 13, 6], [9, 6, 3], [11, 15, 12],
			[15, 11, 13], [15, 13, 14], [4, 7, 1], [7, 4, 11],
			[7, 11, 12], [6, 0, 3], [0, 6, 4], [0, 4, 1], [2, 3, 0],
			[3, 2, 8], [3, 8, 9], [5, 1, 7], [1, 5, 2], [1, 2, 0],
			[10, 12, 15], [12, 10, 5], [12, 5, 7], [8, 14, 9],
			[14, 8, 10], [14, 10, 15], [13, 11, 4, 6], [2, 5, 10, 8]]
	},
	&Polyhedron{
		name:     'j86'
		vertexes: [[f32(-1.10165), f32(-0.110367), f32(-0.010645)],
			[f32(-0.640942), f32(0.825699), f32(0.365159)],
			[f32(-0.414409), f32(0.468967),
				f32(-0.660083)],
			[f32(-0.324965), f32(-0.634882), f32(-0.603383)],
			[f32(-0.317654), f32(-0.702618), f32(0.503439)],
			[f32(0.143053), f32(0.233445),
				f32(0.879242)],
			[f32(0.402426), f32(0.84303), f32(-0.010043)],
			[f32(0.585642), f32(-0.008843),
				f32(-0.69593)],
			[f32(0.603895), f32(-0.925247), f32(-0.07178)],
			[f32(1.0646), f32(0.010817), f32(0.304023)]]
		faces:    [[7, 3, 2], [2, 1, 6], [2, 3, 0], [2, 0, 1],
			[1, 5, 6], [6, 5, 9], [3, 4, 0], [4, 3, 8], [9, 7, 6],
			[9, 8, 7], [7, 8, 3], [6, 7, 2], [1, 0, 4, 5], [5, 4, 8, 9]]
	},
	&Polyhedron{
		name:     'j87'
		vertexes: [[f32(-0.858193), f32(-0.792464), f32(0.432564)],
			[f32(-0.785643), f32(0.057917), f32(-0.211154)],
			[f32(-0.533044), f32(0.147795),
				f32(0.823687)],
			[f32(-0.229952), f32(0.904287), f32(0.131849)],
			[f32(-0.212337), f32(0.637025),
				f32(-0.903062)],
			[f32(-0.091064), f32(-0.748583), f32(-0.310653)],
			[f32(0.161537), f32(-0.658707), f32(0.724189)],
			[f32(0.482242), f32(-0.169476),
				f32(-1.00256)],
			[f32(0.505859), f32(0.352206), f32(0.676436)],
			[f32(0.693906), f32(0.639069),
				f32(-0.336051)],
			[f32(0.86669), f32(-0.369064), f32(-0.025245)]]
		faces:    [[5, 0, 1], [9, 3, 8], [8, 6, 10], [8, 3, 2],
			[8, 2, 6], [6, 5, 10], [10, 5, 7], [3, 1, 2], [1, 3, 4],
			[7, 9, 10], [7, 4, 9], [9, 4, 3], [10, 9, 8], [6, 0, 5],
			[6, 2, 0], [0, 2, 1], [5, 1, 4, 7]]
	},
	&Polyhedron{
		name:     'j88'
		vertexes: [[f32(-0.710639), f32(-0.297668), f32(-0.15267)],
			[f32(-0.651151), f32(-0.105949), f32(0.829841)],
			[f32(-0.621335), f32(0.64788),
				f32(0.169179)],
			[f32(-0.614162), f32(-1.05242), f32(0.500527)],
			[f32(-0.166396), f32(0.361269),
				f32(-0.677289)],
			[f32(-0.002058), f32(-0.993534), f32(-0.291612)],
			[f32(0.165944), f32(0.471894), f32(0.764865)],
			[f32(0.225836), f32(-0.507426),
				f32(0.555374)],
			[f32(0.279224), f32(1.02049), f32(-0.066987)],
			[f32(0.542185), f32(-0.334598),
				f32(-0.816231)],
			[f32(0.770079), f32(0.151511), f32(0.030755)],
			[f32(0.782476), f32(0.638548),
				f32(-0.845752)]]
		faces:    [[6, 7, 10], [3, 7, 1], [3, 5, 7], [10, 11, 8],
			[10, 9, 11], [1, 7, 6], [6, 10, 8], [2, 4, 0], [11, 4, 8],
			[11, 9, 4], [0, 3, 1], [0, 5, 3], [8, 2, 6], [8, 4, 2],
			[2, 1, 6], [2, 0, 1], [7, 5, 9, 10], [4, 9, 5, 0]]
	},
	&Polyhedron{
		name:     'j89'
		vertexes: [[f32(-0.83117), f32(0.133549), f32(-0.011648)],
			[f32(-0.700039), f32(-0.806136), f32(-0.111242)],
			[f32(-0.631074), f32(-0.403619), f32(0.750934)],
			[f32(-0.576095), f32(-0.225432),
				f32(-0.857931)],
			[f32(-0.446282), f32(0.532211), f32(0.764918)],
			[f32(-0.172487), f32(0.817558),
				f32(-0.103263)],
			[f32(0.082589), f32(0.458576), f32(-0.949546)],
			[f32(0.105206), f32(-0.849768),
				f32(-0.620949)],
			[f32(0.145599), f32(-0.76155), f32(0.32811)], [f32(0.235014), f32(-0.09212), f32(1.0019)],
			[f32(0.469795), f32(0.739577), f32(0.597817)],
			[f32(0.750772), f32(0.700456),
				f32(-0.313032)],
			[f32(0.76389), f32(-0.165759), f32(-0.712564)],
			[f32(0.804283), f32(-0.077541),
				f32(0.236495)]]
		faces:    [[9, 8, 13], [1, 8, 2], [1, 7, 8], [13, 11, 10],
			[13, 12, 11], [2, 8, 9], [9, 13, 10], [12, 6, 11],
			[3, 7, 1], [4, 5, 0], [11, 5, 10], [11, 6, 5], [0, 1, 2],
			[0, 3, 1], [10, 4, 9], [10, 5, 4], [4, 2, 9], [4, 0, 2],
			[8, 7, 12, 13], [3, 6, 12, 7], [5, 6, 3, 0]]
	},
	&Polyhedron{
		name:     'j90'
		vertexes: [[f32(-1.05278), f32(0.264006), f32(0.098264)],
			[f32(-0.753999), f32(-0.411397), f32(0.610751)],
			[f32(-0.732127), f32(-0.483215),
				f32(-0.285043)],
			[f32(-0.599216), f32(0.763406), f32(-0.495842)],
			[f32(-0.413906), f32(0.414477),
				f32(0.712494)],
			[f32(-0.278562), f32(0.016184), f32(-0.879148)],
			[f32(-0.105415), f32(-0.890983),
				f32(0.213994)],
			[f32(0.009423), f32(-0.81027), f32(-0.673913)],
			[f32(0.03966), f32(0.913876),
				f32(0.118388)],
			[f32(0.101994), f32(-0.305887), f32(0.864167)],
			[f32(0.267869), f32(0.713733),
				f32(-0.727747)],
			[f32(0.47671), f32(0.507934), f32(0.790906)],
			[f32(0.590474), f32(-0.124774),
				f32(-0.697516)],
			[f32(0.722293), f32(-0.806255), f32(-0.126296)],
			[f32(0.797883), f32(0.460322),
				f32(-0.047343)],
			[f32(0.929701), f32(-0.221158), f32(0.523878)]]
		faces:    [[13, 6, 7], [9, 15, 11], [12, 13, 7], [15, 14, 11],
			[12, 10, 14], [12, 7, 5], [12, 5, 10], [10, 5, 3],
			[7, 6, 2], [5, 7, 2], [2, 6, 1], [2, 1, 0], [10, 3, 8],
			[10, 8, 14], [8, 11, 14], [8, 4, 11], [11, 4, 9],
			[9, 1, 6], [4, 1, 9], [0, 1, 4], [9, 6, 13, 15], [15, 13, 12, 14],
			[5, 2, 0, 3], [3, 0, 4, 8]]
	},
	&Polyhedron{
		name:     'j91'
		vertexes: [[f32(-0.932446), f32(-0.071511), f32(0.062428)],
			[f32(-0.890073), f32(0.716495), f32(0.434115)],
			[f32(-0.483326), f32(0.038238),
				f32(0.802122)],
			[f32(-0.479875), f32(-0.798287), f32(-0.104525)],
			[f32(-0.363346), f32(-0.08879), f32(-0.598427)],
			[f32(-0.294782), f32(1.18623),
				f32(0.002976)],
			[f32(-0.030753), f32(-0.688537), f32(0.635167)],
			[f32(0.030753), f32(0.688538),
				f32(-0.635171)],
			[f32(0.294779), f32(-1.18623), f32(-0.002974)],
			[f32(0.363347), f32(0.088791),
				f32(0.598425)],
			[f32(0.479874), f32(0.79829), f32(0.104525)],
			[f32(0.483327), f32(-0.038241),
				f32(-0.802125)],
			[f32(0.890072), f32(-0.716499), f32(-0.434115)],
			[f32(0.932449), f32(0.071511),
				f32(-0.062429)]]
		faces:    [[11, 13, 12], [7, 11, 4], [10, 7, 5], [13, 10, 9],
			[3, 8, 6], [4, 3, 0], [2, 1, 0], [9, 2, 6], [13, 11, 7, 10],
			[6, 2, 0, 3], [12, 13, 9, 6, 8], [11, 12, 8, 3, 4],
			[5, 7, 4, 0, 1], [10, 5, 1, 2, 9]]
	},
	&Polyhedron{
		name:     'j92'
		vertexes: [[f32(-0.748928), f32(0.557858), f32(-0.030371)],
			[f32(-0.638635), f32(0.125804), f32(-0.670329)],
			[f32(-0.593696), f32(0.259282),
				f32(0.67329)],
			[f32(-0.427424), f32(0.876636), f32(-0.665507)],
			[f32(-0.373109), f32(-0.604827),
				f32(-0.606627)],
			[f32(-0.32817), f32(-0.471348), f32(0.736992)],
			[f32(-0.217876), f32(-0.903403),
				f32(0.097033)],
			[f32(-0.141658), f32(1.0421), f32(0.041134)],
			[f32(-0.021021), f32(0.094954), f32(1.1767)],
			[f32(0.013575), f32(0.743525), f32(0.744795)],
			[f32(0.036802), f32(0.343022),
				f32(-0.994341)],
			[f32(0.267732), f32(-1.03618), f32(-0.498733)],
			[f32(0.302328), f32(-0.387609),
				f32(-0.93064)],
			[f32(0.443205), f32(-0.438661), f32(0.847867)],
			[f32(0.499183), f32(0.610749),
				f32(0.149029)],
			[f32(0.553499), f32(-0.870715), f32(0.207908)],
			[f32(0.609478), f32(0.178694),
				f32(-0.490931)],
			[f32(0.76471), f32(-0.119883), f32(0.212731)]]
		faces:    [[12, 11, 4], [11, 6, 4], [6, 11, 15], [13, 15, 17],
			[5, 13, 8], [2, 5, 8], [2, 8, 9], [7, 9, 14], [16, 14, 17],
			[3, 0, 7], [3, 1, 0], [1, 3, 10], [12, 10, 16], [6, 15, 13, 5],
			[2, 9, 7, 0], [12, 4, 1, 10], [11, 12, 16, 17, 15],
			[8, 13, 17, 14, 9], [16, 10, 3, 7, 14], [1, 4, 6, 5, 2, 0]]
	},
]
